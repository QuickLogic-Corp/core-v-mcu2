/*****************************************************************
          Vendor       : QuickLogic Corp.
          File Name    : top1.vq
          Author       : QuickLogic Corp.

          Description : Verilog Simulation Netlist file
******************************************************************/

`timescale 1ns / 10ps

module top1vq( CLK, RESET, control_in, events_o, fpgaio_in, fpgaio_oe, fpgaio_out, lint_ADDR, lint_BE, lint_GNT, lint_RDATA, lint_REQ, lint_VALID, lint_WDATA, lint_WEN, lint_clk, m0_coef_powerdn, m0_coef_raddr, m0_coef_rclk, m0_coef_rdata, m0_coef_rmode, m0_coef_waddr, m0_coef_wclk, m0_coef_wdata, m0_coef_wdsel, m0_coef_we, m0_coef_wmode, m0_m0_clk, m0_m0_clken, m0_m0_clr, m0_m0_coef_in, m0_m0_csel, m0_m0_dataout, m0_m0_mode, m0_m0_oper_in, m0_m0_osel, m0_m0_outsel, m0_m0_reset, m0_m0_rnd, m0_m0_sat, m0_m0_tc, m0_m1_clk, m0_m1_clken, m0_m1_clr, m0_m1_coef_in, m0_m1_csel, m0_m1_dataout, m0_m1_mode, m0_m1_oper_in, m0_m1_osel, m0_m1_outsel, m0_m1_reset, m0_m1_rnd, m0_m1_sat, m0_m1_tc, m0_oper0_powerdn, m0_oper0_raddr, m0_oper0_rclk, m0_oper0_rdata, m0_oper0_rmode, m0_oper0_waddr, m0_oper0_wclk, m0_oper0_wdata, m0_oper0_wdsel, m0_oper0_we, m0_oper0_wmode, m0_oper1_powerdn, m0_oper1_raddr, m0_oper1_rclk, m0_oper1_rdata, m0_oper1_rmode, m0_oper1_waddr, m0_oper1_wclk, m0_oper1_wdata, m0_oper1_wdsel, m0_oper1_we, m0_oper1_wmode, m1_coef_powerdn, m1_coef_raddr, m1_coef_rclk, m1_coef_rdata, m1_coef_rmode, m1_coef_waddr, m1_coef_wclk, m1_coef_wdata, m1_coef_wdsel, m1_coef_we, m1_coef_wmode, m1_m0_clk, m1_m0_clken, m1_m0_clr, m1_m0_coef_in, m1_m0_csel, m1_m0_dataout, m1_m0_mode, m1_m0_oper_in, m1_m0_osel, m1_m0_outsel, m1_m0_reset, m1_m0_rnd, m1_m0_sat, m1_m0_tc, m1_m1_clk, m1_m1_clken, m1_m1_clr, m1_m1_coef_in, m1_m1_csel, m1_m1_dataout, m1_m1_mode, m1_m1_oper_in, m1_m1_osel, m1_m1_outsel, m1_m1_reset, m1_m1_rnd, m1_m1_sat, m1_m1_tc, m1_oper0_powerdn, m1_oper0_raddr, m1_oper0_rclk, m1_oper0_rdata, m1_oper0_rmode, m1_oper0_waddr, m1_oper0_wclk, m1_oper0_wdata, m1_oper0_wdsel, m1_oper0_we, m1_oper0_wmode, m1_oper1_powerdn, m1_oper1_raddr, m1_oper1_rclk, m1_oper1_rdata, m1_oper1_rmode, m1_oper1_waddr, m1_oper1_wclk, m1_oper1_wdata, m1_oper1_wdsel, m1_oper1_we, m1_oper1_wmode, status_out, tcdm_addr_p0, tcdm_addr_p1, tcdm_addr_p2, tcdm_addr_p3, tcdm_be_p0, tcdm_be_p1, tcdm_be_p2, tcdm_be_p3, tcdm_clk_p0, tcdm_clk_p1, tcdm_clk_p2, tcdm_clk_p3, tcdm_gnt_p0, tcdm_gnt_p1, tcdm_gnt_p2, tcdm_gnt_p3, tcdm_rdata_p0, tcdm_rdata_p1, tcdm_rdata_p2, tcdm_rdata_p3, tcdm_req_p0, tcdm_req_p1, tcdm_req_p2, tcdm_req_p3, tcdm_valid_p0, tcdm_valid_p1, tcdm_valid_p2, tcdm_valid_p3, tcdm_wdata_p0, tcdm_wdata_p1, tcdm_wdata_p2, tcdm_wdata_p3, tcdm_wen_p0, tcdm_wen_p1, tcdm_wen_p2, tcdm_wen_p3, version);
input [5:0] CLK;
input [3:0] RESET;
input [31:0] control_in;
output [15:0] events_o;
input [79:0] fpgaio_in;
output [79:0] fpgaio_oe;
output [79:0] fpgaio_out;
input [19:0] lint_ADDR;
input [3:0] lint_BE;
output lint_GNT;
output [31:0] lint_RDATA;
input lint_REQ;
output lint_VALID;
input [31:0] lint_WDATA;
input lint_WEN;
output lint_clk;
output m0_coef_powerdn;
output [11:0] m0_coef_raddr;
output m0_coef_rclk;
input [31:0] m0_coef_rdata;
output [1:0] m0_coef_rmode;
output [11:0] m0_coef_waddr;
output m0_coef_wclk;
output [31:0] m0_coef_wdata;
output m0_coef_wdsel;
output m0_coef_we;
output [1:0] m0_coef_wmode;
output m0_m0_clk;
output m0_m0_clken;
output m0_m0_clr;
output [31:0] m0_m0_coef_in;
output m0_m0_csel;
input [31:0] m0_m0_dataout;
output [1:0] m0_m0_mode;
output [31:0] m0_m0_oper_in;
output m0_m0_osel;
output [5:0] m0_m0_outsel;
output m0_m0_reset;
output m0_m0_rnd;
output m0_m0_sat;
output m0_m0_tc;
output m0_m1_clk;
output m0_m1_clken;
output m0_m1_clr;
output [31:0] m0_m1_coef_in;
output m0_m1_csel;
input [31:0] m0_m1_dataout;
output [1:0] m0_m1_mode;
output [31:0] m0_m1_oper_in;
output m0_m1_osel;
output [5:0] m0_m1_outsel;
output m0_m1_reset;
output m0_m1_rnd;
output m0_m1_sat;
output m0_m1_tc;
output m0_oper0_powerdn;
output [11:0] m0_oper0_raddr;
output m0_oper0_rclk;
input [31:0] m0_oper0_rdata;
output [1:0] m0_oper0_rmode;
output [11:0] m0_oper0_waddr;
output m0_oper0_wclk;
output [31:0] m0_oper0_wdata;
output m0_oper0_wdsel;
output m0_oper0_we;
output [1:0] m0_oper0_wmode;
output m0_oper1_powerdn;
output [11:0] m0_oper1_raddr;
output m0_oper1_rclk;
input [31:0] m0_oper1_rdata;
output [1:0] m0_oper1_rmode;
output [11:0] m0_oper1_waddr;
output m0_oper1_wclk;
output [31:0] m0_oper1_wdata;
output m0_oper1_wdsel;
output m0_oper1_we;
output [1:0] m0_oper1_wmode;
output m1_coef_powerdn;
output [11:0] m1_coef_raddr;
output m1_coef_rclk;
input [31:0] m1_coef_rdata;
output [1:0] m1_coef_rmode;
output [11:0] m1_coef_waddr;
output m1_coef_wclk;
output [31:0] m1_coef_wdata;
output m1_coef_wdsel;
output m1_coef_we;
output [1:0] m1_coef_wmode;
output m1_m0_clk;
output m1_m0_clken;
output m1_m0_clr;
output [31:0] m1_m0_coef_in;
output m1_m0_csel;
input [31:0] m1_m0_dataout;
output [1:0] m1_m0_mode;
output [31:0] m1_m0_oper_in;
output m1_m0_osel;
output [5:0] m1_m0_outsel;
output m1_m0_reset;
output m1_m0_rnd;
output m1_m0_sat;
output m1_m0_tc;
output m1_m1_clk;
output m1_m1_clken;
output m1_m1_clr;
output [31:0] m1_m1_coef_in;
output m1_m1_csel;
input [31:0] m1_m1_dataout;
output [1:0] m1_m1_mode;
output [31:0] m1_m1_oper_in;
output m1_m1_osel;
output [5:0] m1_m1_outsel;
output m1_m1_reset;
output m1_m1_rnd;
output m1_m1_sat;
output m1_m1_tc;
output m1_oper0_powerdn;
output [11:0] m1_oper0_raddr;
output m1_oper0_rclk;
input [31:0] m1_oper0_rdata;
output [1:0] m1_oper0_rmode;
output [11:0] m1_oper0_waddr;
output m1_oper0_wclk;
output [31:0] m1_oper0_wdata;
output m1_oper0_wdsel;
output m1_oper0_we;
output [1:0] m1_oper0_wmode;
output m1_oper1_powerdn;
output [11:0] m1_oper1_raddr;
output m1_oper1_rclk;
input [31:0] m1_oper1_rdata;
output [1:0] m1_oper1_rmode;
output [11:0] m1_oper1_waddr;
output m1_oper1_wclk;
output [31:0] m1_oper1_wdata;
output m1_oper1_wdsel;
output m1_oper1_we;
output [1:0] m1_oper1_wmode;
output [31:0] status_out;
output [19:0] tcdm_addr_p0;
output [19:0] tcdm_addr_p1;
output [19:0] tcdm_addr_p2;
output [19:0] tcdm_addr_p3;
output [3:0] tcdm_be_p0;
output [3:0] tcdm_be_p1;
output [3:0] tcdm_be_p2;
output [3:0] tcdm_be_p3;
output tcdm_clk_p0;
output tcdm_clk_p1;
output tcdm_clk_p2;
output tcdm_clk_p3;
input tcdm_gnt_p0;
input tcdm_gnt_p1;
input tcdm_gnt_p2;
input tcdm_gnt_p3;
input [31:0] tcdm_rdata_p0;
input [31:0] tcdm_rdata_p1;
input [31:0] tcdm_rdata_p2;
input [31:0] tcdm_rdata_p3;
output tcdm_req_p0;
output tcdm_req_p1;
output tcdm_req_p2;
output tcdm_req_p3;
input tcdm_valid_p0;
input tcdm_valid_p1;
input tcdm_valid_p2;
input tcdm_valid_p3;
output [31:0] tcdm_wdata_p0;
output [31:0] tcdm_wdata_p1;
output [31:0] tcdm_wdata_p2;
output [31:0] tcdm_wdata_p3;
output tcdm_wen_p0;
output tcdm_wen_p1;
output tcdm_wen_p2;
output tcdm_wen_p3;
output [7:0] version;

supply1 VCC;
supply0 GND;

wire CLK_int_0__CAND0_BLSBL_1_padClk;
wire CLK_int_0__CAND0_BLSBL_2_padClk;
wire CLK_int_0__CAND0_BLSBL_3_padClk;
wire CLK_int_0__CAND0_BLSBL_4_padClk;
wire CLK_int_0__CAND0_BLSBL_5_padClk;
wire CLK_int_0__CAND0_BLSBL_6_padClk;
wire CLK_int_0__CAND0_BLSBL_7_padClk;
wire CLK_int_0__CAND0_BLSBL_8_padClk;
wire CLK_int_0__CAND0_BLSBR_10_padClk;
wire CLK_int_0__CAND0_BLSBR_11_padClk;
wire CLK_int_0__CAND0_BLSBR_12_padClk;
wire CLK_int_0__CAND0_BLSBR_13_padClk;
wire CLK_int_0__CAND0_BLSBR_14_padClk;
wire CLK_int_0__CAND0_BLSBR_15_padClk;
wire CLK_int_0__CAND0_BLSBR_16_padClk;
wire CLK_int_0__CAND0_BLSBR_9_padClk;
wire CLK_int_0__CAND0_BLSTL_1_padClk;
wire CLK_int_0__CAND0_BLSTL_2_padClk;
wire CLK_int_0__CAND0_BLSTL_3_padClk;
wire CLK_int_0__CAND0_BLSTL_4_padClk;
wire CLK_int_0__CAND0_BLSTL_5_padClk;
wire CLK_int_0__CAND0_BLSTL_6_padClk;
wire CLK_int_0__CAND0_BLSTL_7_padClk;
wire CLK_int_0__CAND0_BLSTL_8_padClk;
wire CLK_int_0__CAND0_BLSTR_10_padClk;
wire CLK_int_0__CAND0_BLSTR_11_padClk;
wire CLK_int_0__CAND0_BLSTR_12_padClk;
wire CLK_int_0__CAND0_BLSTR_13_padClk;
wire CLK_int_0__CAND0_BLSTR_14_padClk;
wire CLK_int_0__CAND0_BLSTR_15_padClk;
wire CLK_int_0__CAND0_BLSTR_9_padClk;
wire CLK_int_0__CAND0_BRSBL_19_padClk;
wire CLK_int_0__CAND0_BRSBL_24_padClk;
wire CLK_int_0__CAND0_BRSBR_25_padClk;
wire CLK_int_0__CAND0_BRSBR_26_padClk;
wire CLK_int_0__CAND0_BRSBR_27_padClk;
wire CLK_int_0__CAND0_BRSBR_28_padClk;
wire CLK_int_0__CAND0_BRSBR_29_padClk;
wire CLK_int_0__CAND0_BRSBR_30_padClk;
wire CLK_int_0__CAND0_BRSBR_31_padClk;
wire CLK_int_0__CAND0_BRSBR_32_padClk;
wire CLK_int_0__CAND0_BRSTL_19_padClk;
wire CLK_int_0__CAND0_BRSTL_20_padClk;
wire CLK_int_0__CAND0_BRSTL_21_padClk;
wire CLK_int_0__CAND0_BRSTR_29_padClk;
wire CLK_int_0__CAND0_BRSTR_30_padClk;
wire CLK_int_0__CAND0_BRSTR_31_padClk;
wire CLK_int_0__CAND0_BRSTR_32_padClk;
wire CLK_int_0__CAND0_BRSTR_33_padClk;
wire CLK_int_0__CAND0_TLSBL_0_padClk;
wire CLK_int_0__CAND0_TLSBL_1_padClk;
wire CLK_int_0__CAND0_TLSBL_3_padClk;
wire CLK_int_0__CAND0_TLSBL_4_padClk;
wire CLK_int_0__CAND0_TLSBL_5_padClk;
wire CLK_int_0__CAND0_TLSBL_6_padClk;
wire CLK_int_0__CAND0_TLSBL_7_padClk;
wire CLK_int_0__CAND0_TLSBL_8_padClk;
wire CLK_int_0__CAND0_TLSBR_10_padClk;
wire CLK_int_0__CAND0_TLSBR_11_padClk;
wire CLK_int_0__CAND0_TLSBR_12_padClk;
wire CLK_int_0__CAND0_TLSBR_13_padClk;
wire CLK_int_0__CAND0_TLSBR_14_padClk;
wire CLK_int_0__CAND0_TLSBR_15_padClk;
wire CLK_int_0__CAND0_TLSBR_16_padClk;
wire CLK_int_0__CAND0_TLSBR_9_padClk;
wire CLK_int_0__CAND0_TLSTL_1_padClk;
wire CLK_int_0__CAND0_TLSTL_2_padClk;
wire CLK_int_0__CAND0_TLSTL_3_padClk;
wire CLK_int_0__CAND0_TLSTL_4_padClk;
wire CLK_int_0__CAND0_TLSTL_5_padClk;
wire CLK_int_0__CAND0_TLSTL_6_padClk;
wire CLK_int_0__CAND0_TLSTL_7_padClk;
wire CLK_int_0__CAND0_TLSTR_10_padClk;
wire CLK_int_0__CAND0_TLSTR_11_padClk;
wire CLK_int_0__CAND0_TLSTR_12_padClk;
wire CLK_int_0__CAND0_TLSTR_13_padClk;
wire CLK_int_0__CAND0_TLSTR_14_padClk;
wire CLK_int_0__CAND0_TLSTR_15_padClk;
wire CLK_int_0__CAND0_TLSTR_16_padClk;
wire CLK_int_0__CAND0_TRSBL_17_padClk;
wire CLK_int_0__CAND0_TRSBL_18_padClk;
wire CLK_int_0__CAND0_TRSBL_19_padClk;
wire CLK_int_0__CAND0_TRSBL_20_padClk;
wire CLK_int_0__CAND0_TRSBL_21_padClk;
wire CLK_int_0__CAND0_TRSBR_29_padClk;
wire CLK_int_0__CAND0_TRSBR_30_padClk;
wire CLK_int_0__CAND0_TRSBR_31_padClk;
wire CLK_int_0__CAND0_TRSBR_32_padClk;
wire CLK_int_0__CAND0_TRSBR_33_padClk;
wire CLK_int_0__CAND0_TRSTL_17_padClk;
wire CLK_int_0__CAND0_TRSTL_19_padClk;
wire CLK_int_0__CAND0_TRSTL_24_padClk;
wire CLK_int_0__CAND0_TRSTR_25_padClk;
wire CLK_int_0__CAND0_TRSTR_26_padClk;
wire CLK_int_0__CAND0_TRSTR_27_padClk;
wire CLK_int_0__CAND0_TRSTR_28_padClk;
wire CLK_int_0__CAND0_TRSTR_29_padClk;
wire CLK_int_0__CAND0_TRSTR_30_padClk;
wire CLK_int_0__CAND0_TRSTR_31_padClk;
wire CLK_int_0__CAND0_TRSTR_32_padClk;
wire CLK_int_0__CAND0_TRSTR_33_padClk;
wire CLK_int_0__GMUX_0_padClk;
wire CLK_int_0__QMUX_BL0_padClk;
wire CLK_int_0__QMUX_BR0_padClk;
wire CLK_int_0__QMUX_TL0_padClk;
wire CLK_int_0__QMUX_TR0_padClk;
wire CLK_int_0__SQMUX_BLSBL0_padClk;
wire CLK_int_0__SQMUX_BLSBR0_padClk;
wire CLK_int_0__SQMUX_BLSTL0_padClk;
wire CLK_int_0__SQMUX_BLSTR0_padClk;
wire CLK_int_0__SQMUX_BRSBL0_padClk;
wire CLK_int_0__SQMUX_BRSBR0_padClk;
wire CLK_int_0__SQMUX_BRSTL0_padClk;
wire CLK_int_0__SQMUX_BRSTR0_padClk;
wire CLK_int_0__SQMUX_TLSBL0_padClk;
wire CLK_int_0__SQMUX_TLSBR0_padClk;
wire CLK_int_0__SQMUX_TLSTL0_padClk;
wire CLK_int_0__SQMUX_TLSTR0_padClk;
wire CLK_int_0__SQMUX_TRSBL0_padClk;
wire CLK_int_0__SQMUX_TRSBR0_padClk;
wire CLK_int_0__SQMUX_TRSTL0_padClk;
wire CLK_int_0__SQMUX_TRSTR0_padClk;
wire CLK_int_1__CAND1_TLSBL_8_padClk;
wire CLK_int_1__GMUX_1_padClk;
wire CLK_int_1__QMUX_TL1_padClk;
wire CLK_int_1__SQMUX_TLSBL1_padClk;
wire CLK_int_2__CAND2_TLSBR_9_padClk;
wire CLK_int_2__GMUX_2_padClk;
wire CLK_int_2__QMUX_TL2_padClk;
wire CLK_int_2__SQMUX_TLSBR2_padClk;
wire CLK_int_3__CAND3_TLSBL_5_padClk;
wire CLK_int_3__GMUX_3_padClk;
wire CLK_int_3__QMUX_TL3_padClk;
wire CLK_int_3__SQMUX_TLSBL3_padClk;
wire CLK_int_4__CAND4_TLSBL_7_padClk;
wire CLK_int_4__GMUX_4_padClk;
wire CLK_int_4__QMUX_TL4_padClk;
wire CLK_int_4__SQMUX_TLSBL4_padClk;
wire CLK_int_5__CAND5_TLSBR_9_padClk;
wire CLK_int_5__GMUX_5_padClk;
wire CLK_int_5__QMUX_TL5_padClk;
wire CLK_int_5__SQMUX_TLSBR5_padClk;
wire NET_0;
wire NET_1;
wire NET_10;
wire NET_100;
wire NET_101;
wire NET_102;
wire NET_103;
wire NET_104;
wire NET_105;
wire NET_106;
wire NET_107;
wire NET_108;
wire NET_109;
wire NET_11;
wire NET_110;
wire NET_110_CAND3_TLSBR_13_tpGCLKBUF;
wire NET_110_CAND3_TLSBR_14_tpGCLKBUF;
wire NET_110_CAND3_TLSBR_15_tpGCLKBUF;
wire NET_110_CAND3_TLSBR_16_tpGCLKBUF;
wire NET_110_SQMUX_TLSBR3_tpGCLKBUF;
wire NET_111;
wire NET_112;
wire NET_113;
wire NET_114;
wire NET_115;
wire NET_116;
wire NET_117;
wire NET_118;
wire NET_119;
wire NET_12;
wire NET_120;
wire NET_121;
wire NET_122;
wire NET_123;
wire NET_124;
wire NET_125;
wire NET_125_CAND4_TLSBR_13_tpGCLKBUF;
wire NET_125_CAND4_TLSBR_14_tpGCLKBUF;
wire NET_125_CAND4_TLSBR_15_tpGCLKBUF;
wire NET_125_CAND4_TLSBR_16_tpGCLKBUF;
wire NET_125_SQMUX_TLSBR4_tpGCLKBUF;
wire NET_126;
wire NET_127;
wire NET_128;
wire NET_129;
wire NET_13;
wire NET_130;
wire NET_131;
wire NET_132;
wire NET_133;
wire NET_134;
wire NET_135;
wire NET_136;
wire NET_137;
wire NET_138;
wire NET_139;
wire NET_14;
wire NET_140;
wire NET_141;
wire NET_142;
wire NET_143;
wire NET_144;
wire NET_145;
wire NET_146;
wire NET_147;
wire NET_148;
wire NET_149;
wire NET_15;
wire NET_150;
wire NET_151;
wire NET_152;
wire NET_153;
wire NET_154;
wire NET_155;
wire NET_156;
wire NET_157;
wire NET_158;
wire NET_159;
wire NET_16;
wire NET_160;
wire NET_161;
wire NET_162;
wire NET_163;
wire NET_164;
wire NET_165;
wire NET_166;
wire NET_167;
wire NET_168;
wire NET_169;
wire NET_17;
wire NET_170;
wire NET_171;
wire NET_172;
wire NET_173;
wire NET_174;
wire NET_175;
wire NET_176;
wire NET_177;
wire NET_178;
wire NET_179;
wire NET_17_CAND2_BLSTR_10_tpGCLKBUF;
wire NET_17_CAND2_BLSTR_11_tpGCLKBUF;
wire NET_17_CAND2_BLSTR_12_tpGCLKBUF;
wire NET_17_CAND2_BLSTR_13_tpGCLKBUF;
wire NET_17_CAND2_BLSTR_14_tpGCLKBUF;
wire NET_17_CAND2_BLSTR_9_tpGCLKBUF;
wire NET_17_SQMUX_BLSTR2_tpGCLKBUF;
wire NET_18;
wire NET_180;
wire NET_181;
wire NET_182;
wire NET_183;
wire NET_184;
wire NET_185;
wire NET_186;
wire NET_187;
wire NET_188;
wire NET_189;
wire NET_18_CAND4_BLSTR_10_tpGCLKBUF;
wire NET_18_CAND4_BLSTR_11_tpGCLKBUF;
wire NET_18_CAND4_BLSTR_9_tpGCLKBUF;
wire NET_18_SQMUX_BLSTR4_tpGCLKBUF;
wire NET_19;
wire NET_190;
wire NET_191;
wire NET_192;
wire NET_193;
wire NET_194;
wire NET_195;
wire NET_196;
wire NET_197;
wire NET_198;
wire NET_199;
wire NET_2;
wire NET_20;
wire NET_200;
wire NET_201;
wire NET_202;
wire NET_203;
wire NET_204;
wire NET_205;
wire NET_206;
wire NET_207;
wire NET_208;
wire NET_209;
wire NET_21;
wire NET_210;
wire NET_211;
wire NET_212;
wire NET_213;
wire NET_214;
wire NET_215;
wire NET_216;
wire NET_217;
wire NET_218;
wire NET_219;
wire NET_22;
wire NET_220;
wire NET_221;
wire NET_222;
wire NET_223;
wire NET_224;
wire NET_225;
wire NET_226;
wire NET_227;
wire NET_228;
wire NET_229;
wire NET_23;
wire NET_230;
wire NET_231;
wire NET_232;
wire NET_233;
wire NET_234;
wire NET_235;
wire NET_236;
wire NET_237;
wire NET_238;
wire NET_239;
wire NET_24;
wire NET_240;
wire NET_241;
wire NET_242;
wire NET_243;
wire NET_244;
wire NET_245;
wire NET_246;
wire NET_247;
wire NET_248;
wire NET_249;
wire NET_25;
wire NET_250;
wire NET_251;
wire NET_252;
wire NET_253;
wire NET_254;
wire NET_255;
wire NET_256;
wire NET_257;
wire NET_258;
wire NET_259;
wire NET_26;
wire NET_260;
wire NET_261;
wire NET_262;
wire NET_263;
wire NET_264;
wire NET_265;
wire NET_266;
wire NET_267;
wire NET_268;
wire NET_269;
wire NET_27;
wire NET_270;
wire NET_271;
wire NET_272;
wire NET_273;
wire NET_274;
wire NET_275;
wire NET_276;
wire NET_277;
wire NET_278;
wire NET_279;
wire NET_28;
wire NET_280;
wire NET_281;
wire NET_282;
wire NET_283;
wire NET_284;
wire NET_285;
wire NET_286;
wire NET_287;
wire NET_288;
wire NET_289;
wire NET_28_CAND5_BLSTR_12_tpGCLKBUF;
wire NET_28_CAND5_BLSTR_13_tpGCLKBUF;
wire NET_28_CAND5_BLSTR_14_tpGCLKBUF;
wire NET_28_CAND5_BLSTR_9_tpGCLKBUF;
wire NET_28_SQMUX_BLSTR5_tpGCLKBUF;
wire NET_29;
wire NET_290;
wire NET_291;
wire NET_292;
wire NET_293;
wire NET_294;
wire NET_295;
wire NET_296;
wire NET_297;
wire NET_298;
wire NET_299;
wire NET_29_CAND4_BLSTL_2_tpGCLKBUF;
wire NET_29_CAND4_BLSTL_7_tpGCLKBUF;
wire NET_29_CAND4_BLSTL_8_tpGCLKBUF;
wire NET_29_SQMUX_BLSTL4_tpGCLKBUF;
wire NET_3;
wire NET_30;
wire NET_300;
wire NET_301;
wire NET_302;
wire NET_303;
wire NET_304;
wire NET_305;
wire NET_306;
wire NET_307;
wire NET_308;
wire NET_309;
wire NET_31;
wire NET_310;
wire NET_311;
wire NET_312;
wire NET_313;
wire NET_314;
wire NET_315;
wire NET_316;
wire NET_317;
wire NET_318;
wire NET_319;
wire NET_32;
wire NET_320;
wire NET_321;
wire NET_322;
wire NET_323;
wire NET_324;
wire NET_325;
wire NET_326;
wire NET_327;
wire NET_328;
wire NET_329;
wire NET_33;
wire NET_330;
wire NET_331;
wire NET_332;
wire NET_333;
wire NET_334;
wire NET_335;
wire NET_336;
wire NET_337;
wire NET_338;
wire NET_339;
wire NET_34;
wire NET_340;
wire NET_341;
wire NET_342;
wire NET_343;
wire NET_344;
wire NET_345;
wire NET_346;
wire NET_347;
wire NET_348;
wire NET_349;
wire NET_35;
wire NET_350;
wire NET_351;
wire NET_352;
wire NET_353;
wire NET_354;
wire NET_355;
wire NET_356;
wire NET_357;
wire NET_358;
wire NET_359;
wire NET_36;
wire NET_360;
wire NET_361;
wire NET_362;
wire NET_363;
wire NET_364;
wire NET_365;
wire NET_366;
wire NET_367;
wire NET_368;
wire NET_369;
wire NET_37;
wire NET_370;
wire NET_371;
wire NET_372;
wire NET_373;
wire NET_374;
wire NET_375;
wire NET_376;
wire NET_377;
wire NET_378;
wire NET_379;
wire NET_38;
wire NET_380;
wire NET_381;
wire NET_382;
wire NET_383;
wire NET_384;
wire NET_385;
wire NET_386;
wire NET_387;
wire NET_388;
wire NET_389;
wire NET_39;
wire NET_390;
wire NET_391;
wire NET_392;
wire NET_393;
wire NET_394;
wire NET_395;
wire NET_396;
wire NET_397;
wire NET_398;
wire NET_399;
wire NET_4;
wire NET_40;
wire NET_400;
wire NET_401;
wire NET_402;
wire NET_403;
wire NET_404;
wire NET_405;
wire NET_406;
wire NET_407;
wire NET_408;
wire NET_409;
wire NET_41;
wire NET_410;
wire NET_411;
wire NET_412;
wire NET_413;
wire NET_414;
wire NET_415;
wire NET_416;
wire NET_417;
wire NET_418;
wire NET_419;
wire NET_41_CAND4_TLSTR_10_tpGCLKBUF;
wire NET_41_CAND4_TLSTR_11_tpGCLKBUF;
wire NET_41_CAND4_TLSTR_13_tpGCLKBUF;
wire NET_41_CAND4_TLSTR_14_tpGCLKBUF;
wire NET_41_CAND4_TLSTR_15_tpGCLKBUF;
wire NET_41_CAND4_TLSTR_16_tpGCLKBUF;
wire NET_41_SQMUX_TLSTR4_tpGCLKBUF;
wire NET_42;
wire NET_420;
wire NET_421;
wire NET_422;
wire NET_423;
wire NET_424;
wire NET_425;
wire NET_426;
wire NET_427;
wire NET_428;
wire NET_429;
wire NET_43;
wire NET_430;
wire NET_431;
wire NET_432;
wire NET_433;
wire NET_434;
wire NET_435;
wire NET_436;
wire NET_437;
wire NET_438;
wire NET_439;
wire NET_43_CAND3_BLSBR_10_tpGCLKBUF;
wire NET_43_CAND3_BLSBR_11_tpGCLKBUF;
wire NET_43_CAND3_BLSBR_12_tpGCLKBUF;
wire NET_43_CAND3_BLSBR_13_tpGCLKBUF;
wire NET_43_CAND3_BLSBR_14_tpGCLKBUF;
wire NET_43_CAND3_BLSBR_15_tpGCLKBUF;
wire NET_43_CAND3_BLSBR_9_tpGCLKBUF;
wire NET_43_SQMUX_BLSBR3_tpGCLKBUF;
wire NET_44;
wire NET_440;
wire NET_441;
wire NET_442;
wire NET_443;
wire NET_444;
wire NET_445;
wire NET_446;
wire NET_447;
wire NET_448;
wire NET_449;
wire NET_44_CAND4_BLSBR_10_tpGCLKBUF;
wire NET_44_CAND4_BLSBR_11_tpGCLKBUF;
wire NET_44_CAND4_BLSBR_12_tpGCLKBUF;
wire NET_44_CAND4_BLSBR_13_tpGCLKBUF;
wire NET_44_CAND4_BLSBR_14_tpGCLKBUF;
wire NET_44_CAND4_BLSBR_15_tpGCLKBUF;
wire NET_44_SQMUX_BLSBR4_tpGCLKBUF;
wire NET_45;
wire NET_450;
wire NET_451;
wire NET_452;
wire NET_453;
wire NET_454;
wire NET_455;
wire NET_456;
wire NET_457;
wire NET_458;
wire NET_459;
wire NET_45_CAND5_BLSBR_10_tpGCLKBUF;
wire NET_45_CAND5_BLSBR_11_tpGCLKBUF;
wire NET_45_CAND5_BLSBR_9_tpGCLKBUF;
wire NET_45_CAND5_TLSTR_10_tpGCLKBUF;
wire NET_45_CAND5_TLSTR_11_tpGCLKBUF;
wire NET_45_CAND5_TLSTR_9_tpGCLKBUF;
wire NET_45_SQMUX_BLSBR5_tpGCLKBUF;
wire NET_45_SQMUX_TLSTR5_tpGCLKBUF;
wire NET_46;
wire NET_460;
wire NET_461;
wire NET_462;
wire NET_463;
wire NET_464;
wire NET_465;
wire NET_466;
wire NET_467;
wire NET_468;
wire NET_469;
wire NET_46_CAND3_TLSTR_10_tpGCLKBUF;
wire NET_46_CAND3_TLSTR_11_tpGCLKBUF;
wire NET_46_CAND3_TLSTR_13_tpGCLKBUF;
wire NET_46_CAND3_TLSTR_14_tpGCLKBUF;
wire NET_46_CAND3_TLSTR_15_tpGCLKBUF;
wire NET_46_CAND3_TLSTR_16_tpGCLKBUF;
wire NET_46_CAND3_TLSTR_9_tpGCLKBUF;
wire NET_46_SQMUX_TLSTR3_tpGCLKBUF;
wire NET_47;
wire NET_470;
wire NET_471;
wire NET_472;
wire NET_473;
wire NET_474;
wire NET_475;
wire NET_476;
wire NET_477;
wire NET_478;
wire NET_479;
wire NET_48;
wire NET_480;
wire NET_481;
wire NET_482;
wire NET_483;
wire NET_484;
wire NET_485;
wire NET_486;
wire NET_487;
wire NET_488;
wire NET_489;
wire NET_49;
wire NET_490;
wire NET_491;
wire NET_492;
wire NET_493;
wire NET_494;
wire NET_495;
wire NET_496;
wire NET_497;
wire NET_498;
wire NET_499;
wire NET_49_CAND2_BRSTL_19_tpGCLKBUF;
wire NET_49_CAND2_BRSTL_20_tpGCLKBUF;
wire NET_49_CAND2_BRSTL_21_tpGCLKBUF;
wire NET_49_SQMUX_BRSTL2_tpGCLKBUF;
wire NET_5;
wire NET_50;
wire NET_500;
wire NET_501;
wire NET_502;
wire NET_503;
wire NET_504;
wire NET_505;
wire NET_506;
wire NET_507;
wire NET_508;
wire NET_509;
wire NET_50_CAND4_TRSBL_17_tpGCLKBUF;
wire NET_50_CAND4_TRSBL_19_tpGCLKBUF;
wire NET_50_CAND4_TRSBL_20_tpGCLKBUF;
wire NET_50_CAND4_TRSBL_21_tpGCLKBUF;
wire NET_50_SQMUX_TRSBL4_tpGCLKBUF;
wire NET_51;
wire NET_510;
wire NET_511;
wire NET_512;
wire NET_513;
wire NET_514;
wire NET_515;
wire NET_516;
wire NET_517;
wire NET_518;
wire NET_519;
wire NET_52;
wire NET_520;
wire NET_521;
wire NET_522;
wire NET_523;
wire NET_524;
wire NET_525;
wire NET_526;
wire NET_527;
wire NET_528;
wire NET_529;
wire NET_52_CAND2_TRSBL_18_tpGCLKBUF;
wire NET_52_CAND2_TRSBL_19_tpGCLKBUF;
wire NET_52_CAND2_TRSBL_20_tpGCLKBUF;
wire NET_52_CAND2_TRSBL_21_tpGCLKBUF;
wire NET_52_SQMUX_TRSBL2_tpGCLKBUF;
wire NET_53;
wire NET_530;
wire NET_531;
wire NET_532;
wire NET_533;
wire NET_534;
wire NET_535;
wire NET_536;
wire NET_537;
wire NET_538;
wire NET_539;
wire NET_54;
wire NET_540;
wire NET_541;
wire NET_542;
wire NET_543;
wire NET_544;
wire NET_545;
wire NET_546;
wire NET_547;
wire NET_548;
wire NET_549;
wire NET_55;
wire NET_550;
wire NET_551;
wire NET_552;
wire NET_553;
wire NET_554;
wire NET_555;
wire NET_556;
wire NET_557;
wire NET_558;
wire NET_559;
wire NET_56;
wire NET_560;
wire NET_561;
wire NET_562;
wire NET_563;
wire NET_564;
wire NET_565;
wire NET_566;
wire NET_567;
wire NET_568;
wire NET_569;
wire NET_57;
wire NET_570;
wire NET_571;
wire NET_572;
wire NET_573;
wire NET_574;
wire NET_575;
wire NET_576;
wire NET_577;
wire NET_578;
wire NET_579;
wire NET_58;
wire NET_580;
wire NET_581;
wire NET_582;
wire NET_583;
wire NET_584;
wire NET_585;
wire NET_586;
wire NET_587;
wire NET_588;
wire NET_589;
wire NET_59;
wire NET_590;
wire NET_591;
wire NET_592;
wire NET_593;
wire NET_594;
wire NET_595;
wire NET_596;
wire NET_597;
wire NET_598;
wire NET_599;
wire NET_6;
wire NET_60;
wire NET_600;
wire NET_601;
wire NET_602;
wire NET_603;
wire NET_604;
wire NET_605;
wire NET_606;
wire NET_607;
wire NET_608;
wire NET_609;
wire NET_61;
wire NET_610;
wire NET_611;
wire NET_612;
wire NET_613;
wire NET_614;
wire NET_615;
wire NET_616;
wire NET_617;
wire NET_618;
wire NET_619;
wire NET_62;
wire NET_620;
wire NET_621;
wire NET_622;
wire NET_623;
wire NET_624;
wire NET_625;
wire NET_626;
wire NET_627;
wire NET_628;
wire NET_629;
wire NET_63;
wire NET_630;
wire NET_631;
wire NET_632;
wire NET_633;
wire NET_634;
wire NET_635;
wire NET_636;
wire NET_637;
wire NET_638;
wire NET_639;
wire NET_64;
wire NET_640;
wire NET_641;
wire NET_642;
wire NET_643;
wire NET_644;
wire NET_645;
wire NET_646;
wire NET_647;
wire NET_648;
wire NET_649;
wire NET_65;
wire NET_650;
wire NET_651;
wire NET_652;
wire NET_653;
wire NET_654;
wire NET_655;
wire NET_656;
wire NET_657;
wire NET_658;
wire NET_659;
wire NET_66;
wire NET_660;
wire NET_661;
wire NET_662;
wire NET_663;
wire NET_664;
wire NET_665;
wire NET_666;
wire NET_667;
wire NET_668;
wire NET_669;
wire NET_67;
wire NET_670;
wire NET_671;
wire NET_672;
wire NET_673;
wire NET_674;
wire NET_675;
wire NET_676;
wire NET_677;
wire NET_678;
wire NET_679;
wire NET_68;
wire NET_680;
wire NET_681;
wire NET_682;
wire NET_683;
wire NET_684;
wire NET_685;
wire NET_686;
wire NET_687;
wire NET_688;
wire NET_689;
wire NET_69;
wire NET_690;
wire NET_691;
wire NET_692;
wire NET_693;
wire NET_694;
wire NET_695;
wire NET_696;
wire NET_697;
wire NET_698;
wire NET_699;
wire NET_7;
wire NET_70;
wire NET_700;
wire NET_701;
wire NET_702;
wire NET_703;
wire NET_704;
wire NET_705;
wire NET_706;
wire NET_707;
wire NET_708;
wire NET_709;
wire NET_71;
wire NET_710;
wire NET_711;
wire NET_712;
wire NET_713;
wire NET_714;
wire NET_715;
wire NET_716;
wire NET_717;
wire NET_718;
wire NET_719;
wire NET_72;
wire NET_720;
wire NET_721;
wire NET_722;
wire NET_723;
wire NET_724;
wire NET_725;
wire NET_726;
wire NET_727;
wire NET_728;
wire NET_729;
wire NET_73;
wire NET_730;
wire NET_731;
wire NET_732;
wire NET_733;
wire NET_734;
wire NET_735;
wire NET_736;
wire NET_737;
wire NET_738;
wire NET_739;
wire NET_74;
wire NET_740;
wire NET_741;
wire NET_742;
wire NET_743;
wire NET_744;
wire NET_745;
wire NET_746;
wire NET_747;
wire NET_748;
wire NET_749;
wire NET_75;
wire NET_750;
wire NET_751;
wire NET_752;
wire NET_753;
wire NET_754;
wire NET_755;
wire NET_756;
wire NET_757;
wire NET_758;
wire NET_759;
wire NET_76;
wire NET_760;
wire NET_761;
wire NET_762;
wire NET_77;
wire NET_78;
wire NET_79;
wire NET_7_CAND3_BRSTL_19_tpGCLKBUF;
wire NET_7_CAND3_BRSTL_20_tpGCLKBUF;
wire NET_7_CAND3_BRSTL_21_tpGCLKBUF;
wire NET_7_SQMUX_BRSTL3_tpGCLKBUF;
wire NET_8;
wire NET_80;
wire NET_81;
wire NET_82;
wire NET_83;
wire NET_83_CAND3_TRSBL_18_tpGCLKBUF;
wire NET_83_CAND3_TRSBL_19_tpGCLKBUF;
wire NET_83_SQMUX_TRSBL3_tpGCLKBUF;
wire NET_84;
wire NET_85;
wire NET_86;
wire NET_87;
wire NET_88;
wire NET_89;
wire NET_8_CAND5_TLSBL_1_tpGCLKBUF;
wire NET_8_CAND5_TLSBL_2_tpGCLKBUF;
wire NET_8_CAND5_TLSBL_3_tpGCLKBUF;
wire NET_8_CAND5_TLSBL_4_tpGCLKBUF;
wire NET_8_CAND5_TLSBL_7_tpGCLKBUF;
wire NET_8_CAND5_TLSBL_8_tpGCLKBUF;
wire NET_8_SQMUX_TLSBL5_tpGCLKBUF;
wire NET_9;
wire NET_90;
wire NET_91;
wire NET_92;
wire NET_93;
wire NET_94;
wire NET_94_CAND3_BLSTL_5_tpGCLKBUF;
wire NET_94_CAND3_BLSTL_6_tpGCLKBUF;
wire NET_94_CAND3_BLSTL_7_tpGCLKBUF;
wire NET_94_CAND3_BLSTL_8_tpGCLKBUF;
wire NET_94_SQMUX_BLSTL3_tpGCLKBUF;
wire NET_95;
wire NET_96;
wire NET_97;
wire NET_98;
wire NET_99;
wire lint_ADDR_int_11__CAND5_TLSTL_4_tpGCLKBUF;
wire lint_ADDR_int_11__CAND5_TLSTL_5_tpGCLKBUF;
wire lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF;
wire lint_ADDR_int_11__SQMUX_TLSTL5_tpGCLKBUF;
wire lint_GNT;
wire lint_GNT_dup_0;
wire lint_REQ;
wire lint_REQ_int;
wire lint_VALID;
wire lint_VALID_dup_0;
wire lint_WEN;
wire lint_WEN_int;
wire lint_clk;
wire m0_coef_powerdn;
wire m0_coef_rclk;
wire m0_coef_wclk;
wire m0_coef_wdsel;
wire m0_coef_wdsel_dup_0;
wire m0_coef_we;
wire m0_coef_we_dup_0;
wire m0_m0_clk;
wire m0_m0_clken;
wire m0_m0_clken_dup_0;
wire m0_m0_clr;
wire m0_m0_clr_dup_0;
wire m0_m0_csel;
wire m0_m0_csel_dup_0;
wire m0_m0_osel;
wire m0_m0_osel_dup_0;
wire m0_m0_reset;
wire m0_m0_reset_dup_0;
wire m0_m0_rnd;
wire m0_m0_rnd_dup_0;
wire m0_m0_sat;
wire m0_m0_sat_dup_0;
wire m0_m0_tc;
wire m0_m0_tc_dup_0;
wire m0_m1_clk;
wire m0_m1_clken;
wire m0_m1_clken_dup_0;
wire m0_m1_clr;
wire m0_m1_clr_dup_0;
wire m0_m1_csel;
wire m0_m1_csel_dup_0;
wire m0_m1_osel;
wire m0_m1_osel_dup_0;
wire m0_m1_reset;
wire m0_m1_reset_dup_0;
wire m0_m1_rnd;
wire m0_m1_rnd_dup_0;
wire m0_m1_sat;
wire m0_m1_sat_dup_0;
wire m0_m1_tc;
wire m0_m1_tc_dup_0;
wire m0_oper0_powerdn;
wire m0_oper0_rclk;
wire m0_oper0_wclk;
wire m0_oper0_wdsel;
wire m0_oper0_wdsel_dup_0;
wire m0_oper0_we;
wire m0_oper0_we_dup_0;
wire m0_oper1_powerdn;
wire m0_oper1_rclk;
wire m0_oper1_wclk;
wire m0_oper1_wdsel;
wire m0_oper1_wdsel_dup_0;
wire m0_oper1_we;
wire m0_oper1_we_dup_0;
wire m1_coef_powerdn;
wire m1_coef_rclk;
wire m1_coef_wclk;
wire m1_coef_wdsel;
wire m1_coef_we;
wire m1_coef_we_dup_0;
wire m1_m0_clk;
wire m1_m0_clken;
wire m1_m0_clken_dup_0;
wire m1_m0_clr;
wire m1_m0_clr_dup_0;
wire m1_m0_csel;
wire m1_m0_csel_dup_0;
wire m1_m0_osel;
wire m1_m0_osel_dup_0;
wire m1_m0_reset;
wire m1_m0_reset_dup_0;
wire m1_m0_rnd;
wire m1_m0_rnd_dup_0;
wire m1_m0_sat;
wire m1_m0_sat_dup_0;
wire m1_m0_tc;
wire m1_m0_tc_dup_0;
wire m1_m1_clk;
wire m1_m1_clken;
wire m1_m1_clken_dup_0;
wire m1_m1_clr;
wire m1_m1_clr_dup_0;
wire m1_m1_csel;
wire m1_m1_csel_dup_0;
wire m1_m1_osel;
wire m1_m1_osel_dup_0;
wire m1_m1_reset;
wire m1_m1_reset_dup_0;
wire m1_m1_rnd;
wire m1_m1_rnd_dup_0;
wire m1_m1_sat;
wire m1_m1_sat_dup_0;
wire m1_m1_tc;
wire m1_m1_tc_dup_0;
wire m1_oper0_powerdn;
wire m1_oper0_rclk;
wire m1_oper0_wclk;
wire m1_oper0_wdsel;
wire m1_oper0_we;
wire m1_oper0_we_dup_0;
wire m1_oper1_powerdn;
wire m1_oper1_rclk;
wire m1_oper1_wclk;
wire m1_oper1_wdsel;
wire m1_oper1_we;
wire m1_oper1_we_dup_0;
wire not_RESET_0;
wire not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF;
wire not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF;
wire not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF;
wire not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF;
wire not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF;
wire not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF;
wire not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF;
wire not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF;
wire not_RESET_0_QMUX_BL1_tpGCLKBUF;
wire not_RESET_0_QMUX_BR1_tpGCLKBUF;
wire not_RESET_0_QMUX_TR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSBL2_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF;
wire not_RESET_1;
wire not_RESET_2;
wire not_RESET_3;
wire not_apb_fsm_0;
wire not_apb_fsm_1;
wire nx10146z1;
wire nx10146z2;
wire nx10775z1;
wire nx11310z2;
wire nx11311z2;
wire nx11312z2;
wire nx11313z3;
wire nx14650z1;
wire nx15998z1;
wire nx15998z1_CAND2_TLSTR_11_tpGCLKBUF;
wire nx15998z1_CAND2_TLSTR_12_tpGCLKBUF;
wire nx15998z1_CAND2_TLSTR_13_tpGCLKBUF;
wire nx15998z1_CAND2_TLSTR_14_tpGCLKBUF;
wire nx15998z1_SQMUX_TLSTR2_tpGCLKBUF;
wire nx16907z1;
wire nx18281z1;
wire nx18281z1_CAND5_TRSTR_27_tpGCLKBUF;
wire nx18281z1_CAND5_TRSTR_28_tpGCLKBUF;
wire nx18281z1_CAND5_TRSTR_29_tpGCLKBUF;
wire nx18281z1_SQMUX_TRSTR5_tpGCLKBUF;
wire nx19726z1;
wire nx22245z1;
wire nx22245z1_CAND3_BLSBL_2_tpGCLKBUF;
wire nx22245z1_CAND3_BLSBL_3_tpGCLKBUF;
wire nx22245z1_CAND3_BLSBL_4_tpGCLKBUF;
wire nx22245z1_CAND3_BLSBL_5_tpGCLKBUF;
wire nx22245z1_CAND3_BLSBL_6_tpGCLKBUF;
wire nx22245z1_SQMUX_BLSBL3_tpGCLKBUF;
wire nx23147z1;
wire nx2520z1;
wire nx2520z1_CAND2_BRSBR_30_tpGCLKBUF;
wire nx2520z1_CAND2_BRSBR_31_tpGCLKBUF;
wire nx2520z1_CAND2_BRSBR_32_tpGCLKBUF;
wire nx2520z1_CAND2_BRSTR_30_tpGCLKBUF;
wire nx2520z1_CAND2_BRSTR_31_tpGCLKBUF;
wire nx2520z1_CAND2_BRSTR_32_tpGCLKBUF;
wire nx2520z1_QMUX_BR2_tpGCLKBUF;
wire nx2520z1_SQMUX_BRSBR2_tpGCLKBUF;
wire nx2520z1_SQMUX_BRSTR2_tpGCLKBUF;
wire nx25326z1;
wire nx25587z1;
wire nx25587z1_CAND2_TRSTR_25_tpGCLKBUF;
wire nx25587z1_CAND2_TRSTR_26_tpGCLKBUF;
wire nx25587z1_CAND2_TRSTR_27_tpGCLKBUF;
wire nx25587z1_CAND2_TRSTR_28_tpGCLKBUF;
wire nx25587z1_SQMUX_TRSTR2_tpGCLKBUF;
wire nx25788z1;
wire nx25788z1_CAND3_BRSBR_29_tpGCLKBUF;
wire nx25788z1_CAND3_BRSBR_30_tpGCLKBUF;
wire nx25788z1_CAND3_BRSBR_31_tpGCLKBUF;
wire nx25788z1_CAND3_BRSBR_32_tpGCLKBUF;
wire nx25788z1_SQMUX_BRSBR3_tpGCLKBUF;
wire nx28356z1;
wire nx30664z1;
wire nx30664z1_CAND5_BRSBR_25_tpGCLKBUF;
wire nx30664z1_CAND5_BRSBR_26_tpGCLKBUF;
wire nx30664z1_CAND5_BRSBR_27_tpGCLKBUF;
wire nx30664z1_CAND5_BRSBR_28_tpGCLKBUF;
wire nx30664z1_SQMUX_BRSBR5_tpGCLKBUF;
wire nx30923z1;
wire nx30923z1_CAND4_BRSTR_29_tpGCLKBUF;
wire nx30923z1_CAND4_BRSTR_30_tpGCLKBUF;
wire nx30923z1_CAND4_BRSTR_31_tpGCLKBUF;
wire nx30923z1_CAND4_BRSTR_32_tpGCLKBUF;
wire nx30923z1_SQMUX_BRSTR4_tpGCLKBUF;
wire nx32231z1;
wire nx33579z1;
wire nx33579z1_CAND2_BLSBR_11_tpGCLKBUF;
wire nx33579z1_CAND2_BLSBR_12_tpGCLKBUF;
wire nx33579z1_CAND2_BLSBR_13_tpGCLKBUF;
wire nx33579z1_CAND2_BLSBR_14_tpGCLKBUF;
wire nx33579z1_SQMUX_BLSBR2_tpGCLKBUF;
wire nx34006z1;
wire nx34006z1_CAND2_TLSTL_2_tpGCLKBUF;
wire nx34006z1_CAND2_TLSTL_3_tpGCLKBUF;
wire nx34006z1_CAND2_TLSTL_4_tpGCLKBUF;
wire nx34006z1_CAND2_TLSTL_5_tpGCLKBUF;
wire nx34006z1_CAND2_TLSTL_6_tpGCLKBUF;
wire nx34006z1_SQMUX_TLSTL2_tpGCLKBUF;
wire nx34850z1;
wire nx36058z1;
wire nx36058z1_CAND2_TRSBR_29_tpGCLKBUF;
wire nx36058z1_CAND2_TRSBR_30_tpGCLKBUF;
wire nx36058z1_CAND2_TRSBR_31_tpGCLKBUF;
wire nx36058z1_CAND2_TRSBR_32_tpGCLKBUF;
wire nx36058z1_SQMUX_TRSBR2_tpGCLKBUF;
wire nx39840z1;
wire nx39840z1_CAND4_TLSTL_3_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_4_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_5_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_6_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_7_tpGCLKBUF;
wire nx39840z1_SQMUX_TLSTL4_tpGCLKBUF;
wire nx40728z1;
wire nx41193z1;
wire nx41193z1_CAND3_TRSTR_29_tpGCLKBUF;
wire nx41193z1_CAND3_TRSTR_30_tpGCLKBUF;
wire nx41193z1_CAND3_TRSTR_31_tpGCLKBUF;
wire nx41193z1_CAND3_TRSTR_32_tpGCLKBUF;
wire nx41193z1_SQMUX_TRSTR3_tpGCLKBUF;
wire nx44608z1;
wire nx44608z1_CAND3_TLSTL_1_tpGCLKBUF;
wire nx44608z1_CAND3_TLSTL_2_tpGCLKBUF;
wire nx44608z1_CAND3_TLSTL_3_tpGCLKBUF;
wire nx44608z1_CAND3_TLSTL_4_tpGCLKBUF;
wire nx44608z1_CAND3_TLSTL_5_tpGCLKBUF;
wire nx44608z1_CAND3_TLSTL_6_tpGCLKBUF;
wire nx44608z1_SQMUX_TLSTL3_tpGCLKBUF;
wire nx47611z1;
wire nx47611z1_CAND4_TRSTR_30_tpGCLKBUF;
wire nx47611z1_CAND4_TRSTR_31_tpGCLKBUF;
wire nx47611z1_CAND4_TRSTR_32_tpGCLKBUF;
wire nx47611z1_SQMUX_TRSTR4_tpGCLKBUF;
wire nx4939z1;
wire nx4939z1_CAND5_BLSTL_4_tpGCLKBUF;
wire nx4939z1_CAND5_BLSTL_5_tpGCLKBUF;
wire nx4939z1_CAND5_BLSTL_6_tpGCLKBUF;
wire nx4939z1_CAND5_BLSTL_7_tpGCLKBUF;
wire nx4939z1_CAND5_BLSTL_8_tpGCLKBUF;
wire nx4939z1_SQMUX_BLSTL5_tpGCLKBUF;
wire nx49808z64;
wire nx49871z1;
wire nx49871z1_CAND3_BLSTR_10_tpGCLKBUF;
wire nx49871z1_CAND3_BLSTR_11_tpGCLKBUF;
wire nx49871z1_CAND3_BLSTR_12_tpGCLKBUF;
wire nx49871z1_CAND3_BLSTR_13_tpGCLKBUF;
wire nx49871z1_CAND3_BLSTR_14_tpGCLKBUF;
wire nx49871z1_CAND3_BLSTR_9_tpGCLKBUF;
wire nx49871z1_SQMUX_BLSTR3_tpGCLKBUF;
wire nx52746z1;
wire nx52746z1_CAND3_TRSBR_30_tpGCLKBUF;
wire nx52746z1_CAND3_TRSBR_31_tpGCLKBUF;
wire nx52746z1_CAND3_TRSBR_32_tpGCLKBUF;
wire nx52746z1_SQMUX_TRSBR3_tpGCLKBUF;
wire nx53524z1;
wire nx53672z1;
wire nx53672z1_CAND4_BRSBR_27_tpGCLKBUF;
wire nx53672z1_CAND4_BRSBR_28_tpGCLKBUF;
wire nx53672z1_CAND4_BRSBR_29_tpGCLKBUF;
wire nx53672z1_SQMUX_BRSBR4_tpGCLKBUF;
wire nx57881z1;
wire nx57881z1_CAND3_BRSTR_30_tpGCLKBUF;
wire nx57881z1_CAND3_BRSTR_31_tpGCLKBUF;
wire nx57881z1_CAND3_BRSTR_32_tpGCLKBUF;
wire nx57881z1_SQMUX_BRSTR3_tpGCLKBUF;
wire nx58292z1;
wire nx60509z1;
wire nx60831z1;
wire nx60831z1_CAND4_BLSBL_5_tpGCLKBUF;
wire nx60831z1_CAND4_BLSBL_6_tpGCLKBUF;
wire nx60831z1_SQMUX_BLSBL4_tpGCLKBUF;
wire nx65467z1;
wire nx7012z2;
wire nx7012z3;
wire nx8488z1;
wire nx9707z1;
wire nx9707z1_CAND2_BLSBL_1_tpGCLKBUF;
wire nx9707z1_CAND2_BLSBL_2_tpGCLKBUF;
wire nx9707z1_CAND2_BLSBL_3_tpGCLKBUF;
wire nx9707z1_CAND2_BLSBL_5_tpGCLKBUF;
wire nx9707z1_CAND2_BLSBL_6_tpGCLKBUF;
wire nx9707z1_CAND2_BLSTL_1_tpGCLKBUF;
wire nx9707z1_CAND2_BLSTL_2_tpGCLKBUF;
wire nx9707z1_CAND2_BLSTL_3_tpGCLKBUF;
wire nx9707z1_CAND2_BLSTL_4_tpGCLKBUF;
wire nx9707z1_CAND2_BLSTL_5_tpGCLKBUF;
wire nx9707z1_CAND2_BLSTL_6_tpGCLKBUF;
wire nx9707z1_QMUX_BL2_tpGCLKBUF;
wire nx9707z1_SQMUX_BLSBL2_tpGCLKBUF;
wire nx9707z1_SQMUX_BLSTL2_tpGCLKBUF;
wire saved_REQ;
wire tcdm_clk_p0;
wire tcdm_clk_p1;
wire tcdm_clk_p2;
wire tcdm_clk_p3;
wire tcdm_gnt_p0;
wire tcdm_gnt_p0_int;
wire tcdm_gnt_p1;
wire tcdm_gnt_p1_int;
wire tcdm_gnt_p2;
wire tcdm_gnt_p2_int;
wire tcdm_gnt_p3;
wire tcdm_gnt_p3_int;
wire tcdm_req_p0;
wire tcdm_req_p0_dup_0;
wire tcdm_req_p1;
wire tcdm_req_p1_dup_0;
wire tcdm_req_p2;
wire tcdm_req_p2_dup_0;
wire tcdm_req_p3;
wire tcdm_req_p3_dup_0;
wire tcdm_valid_p0;
wire tcdm_valid_p0_int;
wire tcdm_valid_p1;
wire tcdm_valid_p1_int;
wire tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF;
wire tcdm_valid_p1_int_CAND5_TRSBL_19_tpGCLKBUF;
wire tcdm_valid_p1_int_CAND5_TRSBL_20_tpGCLKBUF;
wire tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF;
wire tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF;
wire tcdm_valid_p2;
wire tcdm_valid_p2_int;
wire tcdm_valid_p3;
wire tcdm_valid_p3_int;
wire tcdm_wen_p0;
wire tcdm_wen_p0_dup_0;
wire tcdm_wen_p1;
wire tcdm_wen_p1_dup_0;
wire tcdm_wen_p2;
wire tcdm_wen_p2_dup_0;
wire tcdm_wen_p3;
wire tcdm_wen_p3_dup_0;
wire [5:0] CLK;
wire [5:0] CLK_int;
wire [3:0] RESET;
wire [3:0] RESET_int;
wire [1:0] apb_fsm;
wire [2:0] cnt1;
wire [2:0] cnt2;
wire [2:0] cnt3;
wire [2:0] cnt4;
wire [2:0] cnt5;
wire [31:0] control_in;
wire [31:0] control_in_int;
wire [15:0] events_o;
wire [79:0] fpgaio_in;
wire [79:0] fpgaio_in_int;
wire [79:0] fpgaio_oe;
wire [79:0] fpgaio_oe_dup_0;
wire [79:0] fpgaio_out;
wire [79:0] fpgaio_out_dup_0;
wire [15:0] i_events;
wire [19:0] lint_ADDR;
wire [19:0] lint_ADDR_int;
wire [3:0] lint_BE;
wire [3:0] lint_BE_int;
wire [31:0] lint_RDATA;
wire [31:0] lint_RDATA_dup_0;
wire [31:0] lint_WDATA;
wire [31:0] lint_WDATA_int;
wire [11:0] m0_coef_raddr;
wire [11:0] m0_coef_raddr_dup_0;
wire [31:0] m0_coef_rdata;
wire [31:0] m0_coef_rdata_int;
wire [1:0] m0_coef_rmode;
wire [1:0] m0_coef_rmode_dup_0;
wire [11:0] m0_coef_waddr;
wire [11:0] m0_coef_waddr_dup_0;
wire [31:0] m0_coef_wdata;
wire [31:0] m0_coef_wdata_dup_0;
wire [1:0] m0_coef_wmode;
wire [1:0] m0_coef_wmode_dup_0;
wire [31:0] m0_m0_coef_in;
wire [30:7] m0_m0_control;
wire [31:0] m0_m0_dataout;
wire [31:0] m0_m0_dataout_int;
wire [1:0] m0_m0_mode;
wire [1:0] m0_m0_mode_dup_0;
wire [31:0] m0_m0_oper_in;
wire [5:0] m0_m0_outsel;
wire [5:0] m0_m0_outsel_dup_0;
wire [31:0] m0_m1_coef_in;
wire [30:7] m0_m1_control;
wire [31:0] m0_m1_dataout;
wire [31:0] m0_m1_dataout_int;
wire [1:0] m0_m1_mode;
wire [1:0] m0_m1_mode_dup_0;
wire [31:0] m0_m1_oper_in;
wire [5:0] m0_m1_outsel;
wire [5:0] m0_m1_outsel_dup_0;
wire [11:0] m0_oper0_raddr;
wire [11:0] m0_oper0_raddr_dup_0;
wire [31:0] m0_oper0_rdata;
wire [31:0] m0_oper0_rdata_int;
wire [1:0] m0_oper0_rmode;
wire [1:0] m0_oper0_rmode_dup_0;
wire [11:0] m0_oper0_waddr;
wire [11:0] m0_oper0_waddr_dup_0;
wire [31:0] m0_oper0_wdata;
wire [31:0] m0_oper0_wdata_dup_0;
wire [1:0] m0_oper0_wmode;
wire [1:0] m0_oper0_wmode_dup_0;
wire [11:0] m0_oper1_raddr;
wire [11:0] m0_oper1_raddr_dup_0;
wire [31:0] m0_oper1_rdata;
wire [31:0] m0_oper1_rdata_int;
wire [1:0] m0_oper1_rmode;
wire [1:0] m0_oper1_rmode_dup_0;
wire [11:0] m0_oper1_waddr;
wire [11:0] m0_oper1_waddr_dup_0;
wire [31:0] m0_oper1_wdata;
wire [31:0] m0_oper1_wdata_dup_0;
wire [1:0] m0_oper1_wmode;
wire [1:0] m0_oper1_wmode_dup_0;
wire [31:15] m0_ram_control;
wire [11:0] m1_coef_raddr;
wire [11:0] m1_coef_raddr_dup_0;
wire [31:0] m1_coef_rdata;
wire [31:0] m1_coef_rdata_int;
wire [1:0] m1_coef_rmode;
wire [11:0] m1_coef_waddr;
wire [11:0] m1_coef_waddr_dup_0;
wire [31:0] m1_coef_wdata;
wire [31:0] m1_coef_wdata_dup_0;
wire [1:0] m1_coef_wmode;
wire [31:0] m1_m0_coef_in;
wire [30:7] m1_m0_control;
wire [31:0] m1_m0_dataout;
wire [31:0] m1_m0_dataout_int;
wire [1:0] m1_m0_mode;
wire [1:0] m1_m0_mode_dup_0;
wire [31:0] m1_m0_oper_in;
wire [5:0] m1_m0_outsel;
wire [5:0] m1_m0_outsel_dup_0;
wire [31:0] m1_m1_coef_in;
wire [30:0] m1_m1_control;
wire [31:0] m1_m1_dataout;
wire [31:0] m1_m1_dataout_int;
wire [1:0] m1_m1_mode;
wire [1:0] m1_m1_mode_dup_0;
wire [31:0] m1_m1_oper_in;
wire [5:0] m1_m1_outsel;
wire [11:0] m1_oper0_raddr;
wire [11:0] m1_oper0_raddr_dup_0;
wire [31:0] m1_oper0_rdata;
wire [31:0] m1_oper0_rdata_int;
wire [1:0] m1_oper0_rmode;
wire [11:0] m1_oper0_waddr;
wire [11:0] m1_oper0_waddr_dup_0;
wire [31:0] m1_oper0_wdata;
wire [31:0] m1_oper0_wdata_dup_0;
wire [1:0] m1_oper0_wmode;
wire [11:0] m1_oper1_raddr;
wire [11:0] m1_oper1_raddr_dup_0;
wire [31:0] m1_oper1_rdata;
wire [31:0] m1_oper1_rdata_int;
wire [1:0] m1_oper1_rmode;
wire [11:0] m1_oper1_waddr;
wire [11:0] m1_oper1_waddr_dup_0;
wire [31:0] m1_oper1_wdata;
wire [31:0] m1_oper1_wdata_dup_0;
wire [1:0] m1_oper1_wmode;
wire [31:0] m1_ram_control;
wire [31:0] status_out;
wire [31:0] status_out_dup_0;
wire [19:0] tcdm_addr_p0;
wire [19:0] tcdm_addr_p0_dup_0;
wire [19:0] tcdm_addr_p1;
wire [19:0] tcdm_addr_p1_dup_0;
wire [19:0] tcdm_addr_p2;
wire [19:0] tcdm_addr_p2_dup_0;
wire [19:0] tcdm_addr_p3;
wire [19:0] tcdm_addr_p3_dup_0;
wire [3:0] tcdm_be_p0;
wire [3:0] tcdm_be_p0_dup_0;
wire [3:0] tcdm_be_p1;
wire [3:0] tcdm_be_p1_dup_0;
wire [3:0] tcdm_be_p2;
wire [3:0] tcdm_be_p2_dup_0;
wire [3:0] tcdm_be_p3;
wire [3:0] tcdm_be_p3_dup_0;
wire [31:0] tcdm_rdata_p0;
wire [31:0] tcdm_rdata_p0_int;
wire [31:0] tcdm_rdata_p1;
wire [31:0] tcdm_rdata_p1_int;
wire [31:0] tcdm_rdata_p2;
wire [31:0] tcdm_rdata_p2_int;
wire [31:0] tcdm_rdata_p3;
wire [31:0] tcdm_rdata_p3_int;
wire [31:0] tcdm_result_p0;
wire [31:0] tcdm_result_p1;
wire [31:0] tcdm_result_p2;
wire [31:0] tcdm_result_p3;
wire [31:0] tcdm_wdata_p0;
wire [31:0] tcdm_wdata_p0_dup_0;
wire [31:0] tcdm_wdata_p1;
wire [31:0] tcdm_wdata_p1_dup_0;
wire [31:0] tcdm_wdata_p2;
wire [31:0] tcdm_wdata_p2_dup_0;
wire [31:0] tcdm_wdata_p3;
wire [31:0] tcdm_wdata_p3_dup_0;
wire [7:0] version;

	LOGIC_0 QL_INST_A4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[19]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[20]),.Q3EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A8_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_oe_dup_0[25]),.B0I1(NET_64),.B0I2(NET_30),.B0I3(fpgaio_in_int[25]),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_oe_dup_0[25]),.T0I1(NET_64),.T0I2(NET_30),.T0I3(fpgaio_in_int[25]),.TB0S(NET_8),.C0Z(NET_506),.Q0Z(fpgaio_oe_dup_0[31]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A8_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(NET_30),.B1I1(NET_64),.B1I2(fpgaio_oe_dup_0[27]),.B1I3(fpgaio_in_int[27]),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_oe_dup_0[27]),.T1I1(fpgaio_in_int[27]),.T1I2(NET_30),.T1I3(NET_64),.TB1S(NET_8),.C1Z(NET_542),.Q1Z(fpgaio_oe_dup_0[18]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_A8_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B2I0(fpgaio_oe_dup_0[31]),.B2I1(NET_64),.B2I2(NET_30),.B2I3(fpgaio_in_int[31]),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_oe_dup_0[31]),.T2I1(NET_64),.T2I2(NET_30),.T2I3(fpgaio_in_int[31]),.TB2S(NET_8),.C2Z(NET_613),.Q2Z(fpgaio_oe_dup_0[22]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_A8_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B3I0(NET_30),.B3I1(fpgaio_oe_dup_0[30]),.B3I2(fpgaio_in_int[30]),.B3I3(NET_64),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_in_int[30]),.T3I1(NET_64),.T3I2(NET_30),.T3I3(fpgaio_oe_dup_0[30]),.TB3S(NET_8),.C3Z(NET_595),.Q3Z(fpgaio_oe_dup_0[30]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_A9_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_10),.B0I1(fpgaio_in_int[37]),.B0I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.B0I3(fpgaio_in_int[5]),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(NET_10),.T0I1(fpgaio_in_int[37]),.T0I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T0I3(fpgaio_in_int[5]),.TB0S(NET_64),.C0Z(NET_661),.Q0Z(fpgaio_oe_dup_0[23]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A9_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B1I0(fpgaio_in_int[3]),.B1I1(NET_10),.B1I2(fpgaio_in_int[35]),.B1I3(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_in_int[35]),.T1I1(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T1I2(fpgaio_in_int[3]),.T1I3(NET_10),.TB1S(NET_64),.C1Z(NET_700),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_A9_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_10),.B2I1(fpgaio_in_int[33]),.B2I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.B2I3(fpgaio_in_int[1]),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.T2I0(NET_10),.T2I1(fpgaio_in_int[33]),.T2I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T2I3(fpgaio_in_int[1]),.TB2S(NET_64),.C2Z(NET_53),.Q2Z(fpgaio_oe_dup_0[24]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_A9_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B3I0(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.B3I1(fpgaio_in_int[36]),.B3I2(NET_10),.B3I3(fpgaio_in_int[4]),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.T3I0(NET_10),.T3I1(fpgaio_in_int[4]),.T3I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T3I3(fpgaio_in_int[36]),.TB3S(NET_64),.C3Z(NET_681),.Q3Z(fpgaio_oe_dup_0[29]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_A10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A10_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_10),.B2I1(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.B2I2(fpgaio_in_int[10]),.B2I3(fpgaio_in_int[42]),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.T2I0(NET_10),.T2I1(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T2I2(fpgaio_in_int[10]),.T2I3(fpgaio_in_int[42]),.TB2S(NET_64),.C2Z(NET_189),.Q2Z(fpgaio_oe_dup_0[21]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_A10_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B3I0(fpgaio_in_int[11]),.B3I1(fpgaio_in_int[43]),.B3I2(NET_10),.B3I3(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.T3I0(NET_10),.T3I1(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T3I2(fpgaio_in_int[11]),.T3I3(fpgaio_in_int[43]),.TB3S(NET_64),.C3Z(NET_208),.Q3Z(fpgaio_oe_dup_0[17]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_A11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A11_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.B1I1(NET_10),.B1I2(fpgaio_in_int[13]),.B1I3(fpgaio_in_int[45]),.T1I0(fpgaio_in_int[13]),.T1I1(fpgaio_in_int[45]),.T1I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T1I3(NET_10),.TB1S(NET_64),.C1Z(NET_248),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_A11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(fpgaio_oe_dup_0[29]),.B2I1(fpgaio_oe_dup_0[61]),.B2I2(NET_123),.B2I3(NET_126),.B2Z(NET_576),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A11_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B3I0(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.B3I1(NET_10),.B3I2(fpgaio_in_int[47]),.B3I3(fpgaio_in_int[15]),.T3I0(fpgaio_in_int[47]),.T3I1(fpgaio_in_int[15]),.T3I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T3I3(NET_10),.TB3S(NET_64),.C3Z(NET_306),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_A12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_123),.B0I1(fpgaio_oe_dup_0[55]),.B0I2(NET_126),.B0I3(fpgaio_oe_dup_0[23]),.B0Z(NET_448),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A12_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(fpgaio_oe_dup_0[18]),.T1I1(fpgaio_oe_dup_0[50]),.T1I2(NET_126),.T1I3(NET_123),.C1Z(NET_358),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_A12_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B2I0(fpgaio_oe_dup_0[17]),.B2I1(fpgaio_oe_dup_0[49]),.B2I2(NET_126),.B2I3(NET_123),.T2I0(NET_123),.T2I1(NET_126),.T2I2(fpgaio_oe_dup_0[22]),.T2I3(fpgaio_oe_dup_0[54]),.TB2S(GND),.B2Z(NET_340),.C2Z(NET_430),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_A12_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_123),.T3I1(NET_126),.T3I2(fpgaio_oe_dup_0[60]),.T3I3(fpgaio_oe_dup_0[28]),.C3Z(NET_558),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_A13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(fpgaio_oe_dup_0[21]),.B0I1(NET_123),.B0I2(NET_126),.B0I3(fpgaio_oe_dup_0[53]),.B0Z(NET_412),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A13_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(fpgaio_oe_dup_0[19]),.T1I1(NET_123),.T1I2(fpgaio_oe_dup_0[51]),.T1I3(NET_126),.C1Z(NET_377),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_A13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_126),.B2I1(NET_123),.B2I2(fpgaio_oe_dup_0[56]),.B2I3(fpgaio_oe_dup_0[24]),.B2Z(NET_487),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A13_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(fpgaio_oe_dup_0[26]),.T3I1(NET_123),.T3I2(NET_126),.T3I3(fpgaio_oe_dup_0[58]),.C3Z(NET_522),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_A14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A14_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.B2I1(fpgaio_in_int[9]),.B2I2(NET_10),.B2I3(fpgaio_in_int[41]),.T2I0(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T2I1(fpgaio_in_int[9]),.T2I2(NET_10),.T2I3(fpgaio_in_int[41]),.TB2S(NET_64),.C2Z(NET_166),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_A14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A15_1 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_30),.T1I1(NET_10),.T1I2(lint_ADDR_int[11]),.T1I3(GND),.C1Z(NET_126),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_A15_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_10),.B2I1(fpgaio_in_int[40]),.B2I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.B2I3(fpgaio_in_int[8]),.T2I0(NET_10),.T2I1(fpgaio_in_int[40]),.T2I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T2I3(fpgaio_in_int[8]),.TB2S(NET_64),.C2Z(NET_287),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_A15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A16_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B0I0(fpgaio_in_int[46]),.B0I1(NET_10),.B0I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.B0I3(fpgaio_in_int[14]),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx9707z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_in_int[46]),.T0I1(NET_10),.T0I2(NET_8_CAND5_TLSBL_1_tpGCLKBUF),.T0I3(fpgaio_in_int[14]),.TB0S(NET_64),.C0Z(NET_268),.Q0Z(fpgaio_oe_dup_0[58]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[24]),.Q3EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[56]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A18_1 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T1I0(NET_10),.T1I1(GND),.T1I2(lint_ADDR_int[11]),.T1I3(NET_64),.C1Z(NET_127),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_A18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[53]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A19_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000001),.B0I0(control_in_int[2]),.B0I1(GND),.B0I2(GND),.B0I3(GND),.T0I0(control_in_int[4]),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND),.B0Z(status_out_dup_0[2]),.C0Z(status_out_dup_0[4]),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_A19_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(control_in_int[0]),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND),.C1Z(status_out_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_A19_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000001),.B2I0(control_in_int[1]),.B2I1(GND),.B2I2(GND),.B2I3(GND),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(control_in_int[5]),.TB2S(GND),.B2Z(status_out_dup_0[1]),.C2Z(status_out_dup_0[5]),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_A19_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(GND),.T3I1(GND),.T3I2(control_in_int[3]),.T3I3(GND),.C3Z(status_out_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_A20_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000001),.B0I0(control_in_int[8]),.B0I1(GND),.B0I2(GND),.B0I3(GND),.T0I0(control_in_int[10]),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND),.B0Z(status_out_dup_0[8]),.C0Z(status_out_dup_0[10]),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_A20_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(GND),.T1I1(GND),.T1I2(control_in_int[13]),.T1I3(GND),.TB1S(GND),.C1Z(status_out_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_A20_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000001),.B2I0(control_in_int[6]),.B2I1(GND),.B2I2(GND),.B2I3(GND),.T2I0(control_in_int[9]),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(status_out_dup_0[6]),.C2Z(status_out_dup_0[9]),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_A20_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(GND),.T3I1(GND),.T3I2(control_in_int[11]),.T3I3(GND),.C3Z(status_out_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_A21_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000001),.B0I0(control_in_int[14]),.B0I1(GND),.B0I2(GND),.B0I3(GND),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(control_in_int[28]),.TB0S(GND),.B0Z(status_out_dup_0[14]),.C0Z(status_out_dup_0[28]),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A21_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T1I0(control_in_int[16]),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND),.C1Z(status_out_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_A21_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000001),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(control_in_int[17]),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(control_in_int[15]),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(status_out_dup_0[17]),.C2Z(status_out_dup_0[15]),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_A21_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T3I0(control_in_int[18]),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND),.C3Z(status_out_dup_0[18]),.Q3Z(fpgaio_oe_dup_0[51]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_A22_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000001),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(control_in_int[25]),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T0I0(control_in_int[20]),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND),.B0Z(status_out_dup_0[25]),.C0Z(status_out_dup_0[20]),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A22_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T1I0(control_in_int[21]),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND),.C1Z(status_out_dup_0[21]),.Q1Z(fpgaio_oe_dup_0[60]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_A22_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000001),.B2I0(GND),.B2I1(control_in_int[22]),.B2I2(GND),.B2I3(GND),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(control_in_int[24]),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(status_out_dup_0[22]),.C2Z(status_out_dup_0[24]),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_A22_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T3I0(control_in_int[23]),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND),.C3Z(status_out_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_A23_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T0I0(control_in_int[29]),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND),.C0Z(status_out_dup_0[29]),.Q0Z(fpgaio_oe_dup_0[55]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A23_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(GND),.T1I2(control_in_int[30]),.T1I3(GND),.TB1S(GND),.C1Z(status_out_dup_0[30]),.Q1Z(fpgaio_oe_dup_0[61]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_A23_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(control_in_int[31]),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND),.C2Z(status_out_dup_0[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_A23_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T3I0(control_in_int[27]),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND),.C3Z(status_out_dup_0[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_A24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[17]),.Q0EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[49]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[50]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[54]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A25_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(NET_127),.T0I1(fpgaio_in_int[39]),.T0I2(fpgaio_oe_dup_0[39]),.T0I3(NET_126),.TB0S(GND),.C0Z(NET_476),.Q0Z(fpgaio_oe_dup_0[34]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A25_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.T1I0(NET_126),.T1I1(NET_127),.T1I2(fpgaio_in_int[44]),.T1I3(fpgaio_oe_dup_0[44]),.TB1S(GND),.C1Z(NET_232),.Q1Z(fpgaio_oe_dup_0[32]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_A25_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B2I0(fpgaio_oe_dup_0[34]),.B2I1(NET_127),.B2I2(fpgaio_in_int[34]),.B2I3(NET_126),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.T2I0(NET_127),.T2I1(fpgaio_in_int[38]),.T2I2(fpgaio_oe_dup_0[38]),.T2I3(NET_126),.TB2S(GND),.B2Z(NET_724),.C2Z(NET_642),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_A25_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.T3I0(NET_127),.T3I1(fpgaio_in_int[32]),.T3I2(fpgaio_oe_dup_0[32]),.T3I3(NET_126),.TB3S(GND),.C3Z(NET_122),.Q3Z(fpgaio_oe_dup_0[44]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_A26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[39]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[38]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[20]),.Q3EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[29]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx44608z1_CAND3_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx44608z1_CAND3_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx44608z1_CAND3_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx44608z1_CAND3_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B8_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(NET_64),.B1I1(NET_30),.B1I2(fpgaio_in_int[20]),.B1I3(fpgaio_oe_dup_0[20]),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx44608z1_CAND3_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_in_int[20]),.T1I1(fpgaio_oe_dup_0[20]),.T1I2(NET_64),.T1I3(NET_30),.TB1S(NET_8),.C1Z(NET_396),.Q1Z(fpgaio_oe_dup_0[0]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_B8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B8_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B3I0(fpgaio_in_int[16]),.B3I1(NET_30),.B3I2(fpgaio_oe_dup_0[16]),.B3I3(NET_64),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_oe_dup_0[16]),.T3I1(NET_64),.T3I2(fpgaio_in_int[16]),.T3I3(NET_30),.TB3S(NET_8),.C3Z(NET_323),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_B9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B2I0(NET_8_CAND5_TLSBL_2_tpGCLKBUF),.B2I1(lint_ADDR_int[11]),.B2I2(GND),.B2I3(NET_30),.B2Z(NET_123),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B11_3 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int[6]),.T3I1(lint_ADDR_int[4]),.T3I2(lint_ADDR_int[3]),.T3I3(lint_ADDR_int[5]),.TB3S(GND),.C3Z(NET_64),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_B18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.B0I1(fpgaio_oe_dup_0[62]),.B0I2(fpgaio_in_int[62]),.B0I3(NET_322),.T0I0(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.T0I1(fpgaio_oe_dup_0[62]),.T0I2(fpgaio_in_int[62]),.T0I3(NET_322),.TB0S(NET_595),.C0Z(NET_593),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_B18_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_64),.T1I1(GND),.T1I2(NET_10),.T1I3(GND),.C1Z(NET_322),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_B18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.B2I1(fpgaio_oe_dup_0[57]),.B2I2(NET_322),.B2I3(fpgaio_in_int[57]),.T2I0(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.T2I1(fpgaio_oe_dup_0[57]),.T2I2(NET_322),.T2I3(fpgaio_in_int[57]),.TB2S(NET_506),.C2Z(NET_504),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_B18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_322),.B0I1(fpgaio_in_int[52]),.B0I2(fpgaio_oe_dup_0[52]),.B0I3(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.T0I0(NET_322),.T0I1(fpgaio_in_int[52]),.T0I2(fpgaio_oe_dup_0[52]),.T0I3(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.TB0S(NET_396),.C0Z(NET_394),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_B19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B1I0(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.B1I1(NET_322),.B1I2(fpgaio_oe_dup_0[59]),.B1I3(fpgaio_in_int[59]),.T1I0(fpgaio_oe_dup_0[59]),.T1I1(fpgaio_in_int[59]),.T1I2(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.T1I3(NET_322),.TB1S(NET_542),.C1Z(NET_540),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_B19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_322),.B2I1(fpgaio_oe_dup_0[63]),.B2I2(fpgaio_in_int[63]),.B2I3(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.T2I0(NET_322),.T2I1(fpgaio_oe_dup_0[63]),.T2I2(fpgaio_in_int[63]),.T2I3(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.TB2S(NET_613),.C2Z(NET_611),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_B19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(fpgaio_in_int[48]),.B3I1(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.B3I2(NET_322),.B3I3(fpgaio_oe_dup_0[48]),.T3I0(NET_322),.T3I1(fpgaio_oe_dup_0[48]),.T3I2(fpgaio_in_int[48]),.T3I3(NET_29_CAND4_BLSTL_2_tpGCLKBUF),.TB3S(NET_323),.C3Z(NET_320),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_B20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B20_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(GND),.T1I2(control_in_int[12]),.T1I3(GND),.TB1S(GND),.C1Z(status_out_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_B20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B20_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx9707z1_CAND2_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.T3I0(control_in_int[7]),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND),.C3Z(status_out_dup_0[7]),.Q3Z(fpgaio_oe_dup_0[57]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_B21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B21_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(control_in_int[19]),.TB2S(GND),.C2Z(status_out_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_B21_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(GND),.T3I1(GND),.T3I2(control_in_int[26]),.T3I3(GND),.TB3S(GND),.C3Z(status_out_dup_0[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_B22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx9707z1_CAND2_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[48]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx9707z1_CAND2_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[63]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[30]),.Q2EN(nx9707z1_CAND2_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[62]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx9707z1_CAND2_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[59]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx9707z1_CAND2_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[52]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx9707z1_CAND2_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[37]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[23]),.Q1EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[23]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[28]),.Q0EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[28]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[30]),.Q2EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[30]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[21]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[10]),.Q1EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_waddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[18]),.Q2EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[18]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[8]),.Q1EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[12]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx44608z1_CAND3_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx39840z1_CAND4_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx39840z1_CAND4_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx39840z1_CAND4_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C8_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.T1I0(NET_124),.T1I1(tcdm_rdata_p0_int[7]),.T1I2(fpgaio_oe_dup_0[7]),.T1I3(NET_123),.C1Z(NET_475),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_C8_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[30]),.Q2EN(nx39840z1_CAND4_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.T2I0(NET_124),.T2I1(fpgaio_oe_dup_0[2]),.T2I2(NET_123),.T2I3(tcdm_rdata_p0_int[2]),.TB2S(GND),.C2Z(NET_723),.Q2Z(fpgaio_out_dup_0[30]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_C8_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_oe_dup_0[6]),.T3I1(tcdm_rdata_p0_int[6]),.T3I2(NET_124),.T3I3(NET_123),.C3Z(NET_641),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_C9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdsel_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.Q0Z(m1_m1_control[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C11_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.T2I0(m1_m1_control[21]),.T2I1(fpgaio_in_int[21]),.T2I2(NET_111),.T2I3(NET_129),.TB2S(GND),.C2Z(NET_415),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_C11_3 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[11]),.T3I1(NET_64),.T3I2(NET_8_CAND5_TLSBL_3_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.C3Z(NET_111),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_C12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.Q0Z(m1_m1_control[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C12_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[23]),.T2I1(m1_m1_control[23]),.T2I2(NET_111),.T2I3(NET_129),.TB2S(GND),.C2Z(NET_451),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_C12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C13_0 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.T0I0(NET_475),.T0I1(GND),.T0I2(NET_474),.T0I3(NET_476),.TB0S(GND),.C0Z(NET_457),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_C13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_rmode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_103),.B0I1(fpgaio_out_dup_0[2]),.B0I2(m0_oper0_wmode_dup_0[0]),.B0I3(NET_102),.B0Z(NET_710),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C14_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_103),.T1I1(fpgaio_out_dup_0[0]),.T1I2(m0_oper0_rmode_dup_0[0]),.T1I3(NET_102),.C1Z(NET_90),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_C14_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.T2I0(fpgaio_out_dup_0[12]),.T2I1(m0_oper0_wdsel_dup_0),.T2I2(NET_103),.T2I3(NET_102),.TB2S(GND),.C2Z(NET_218),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_C14_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_723),.T3I1(NET_724),.T3I2(NET_722),.T3I3(GND),.TB3S(GND),.C3Z(NET_705),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_C15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(m1_m1_control[7]),.B0I1(NET_128),.B0I2(NET_129),.B0I3(fpgaio_out_dup_0[71]),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.T0I0(m1_m1_control[7]),.T0I1(NET_128),.T0I2(NET_129),.T0I3(fpgaio_out_dup_0[71]),.TB0S(NET_477),.C0Z(NET_474),.Q0Z(m1_m1_control[2]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_C15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B1I0(NET_129),.B1I1(fpgaio_out_dup_0[70]),.B1I2(m1_m1_tc_dup_0),.B1I3(NET_128),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_tc_dup_0),.T1I1(NET_128),.T1I2(NET_129),.T1I3(fpgaio_out_dup_0[70]),.TB1S(NET_643),.C1Z(NET_640),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_C15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_m1_control[2]),.B2I1(NET_128),.B2I2(NET_129),.B2I3(fpgaio_out_dup_0[66]),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.T2I0(m1_m1_control[2]),.T2I1(NET_128),.T2I2(NET_129),.T2I3(fpgaio_out_dup_0[66]),.TB2S(NET_725),.C2Z(NET_722),.Q2Z(m1_m1_control[7]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_C15_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.T3I0(NET_641),.T3I1(GND),.T3I2(NET_640),.T3I3(NET_642),.TB3S(GND),.C3Z(NET_623),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_C16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[70]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[76]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[71]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[66]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[67]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[64]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[64]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[75]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[71]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[73]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[77]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[78]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[69]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_rmode_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wmode_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx9707z1_CAND2_BLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[41]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx9707z1_CAND2_BLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[42]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx9707z1_CAND2_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[35]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx9707z1_CAND2_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[46]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[18]),.Q2EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[18]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[9]),.Q1EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[9]),.Q2EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_waddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[4]),.Q0EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_waddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[3]),.Q1EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_waddr_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[9]),.Q2EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_waddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[7]),.Q3EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_waddr_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int_11__CAND5_TLSTL_4_tpGCLKBUF),.Q0EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_waddr_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[6]),.Q1EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_waddr_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[8]),.Q2EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_waddr_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[2]),.Q3EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_waddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx44608z1_CAND3_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[9]),.Q1EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000001000000),.B0I0(lint_ADDR_int[5]),.B0I1(lint_ADDR_int[6]),.B0I2(lint_ADDR_int[4]),.B0I3(lint_ADDR_int[3]),.B0Z(NET_30),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D8_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_123),.T1I1(NET_124),.T1I2(fpgaio_oe_dup_0[0]),.T1I3(tcdm_rdata_p0_int[0]),.C1Z(NET_121),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_D8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_123),.B2I1(NET_124),.B2I2(fpgaio_oe_dup_0[12]),.B2I3(tcdm_rdata_p0_int[12]),.B2Z(NET_231),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[26]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D11_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T0I0(NET_111),.T0I1(NET_129),.T0I2(m1_m1_control[29]),.T0I3(fpgaio_in_int[29]),.TB0S(GND),.C0Z(NET_579),.Q0Z(m1_m1_control[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_D11_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T1I0(RESET_int[3]),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND),.C1Z(not_RESET_3),.Q1Z(m1_m1_control[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_D11_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[24]),.T2I1(m1_m1_control[24]),.T2I2(NET_111),.T2I3(NET_129),.TB2S(GND),.C2Z(NET_490),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_D11_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T3I0(NET_111),.T3I1(m1_m1_control[28]),.T3I2(fpgaio_in_int[28]),.T3I3(NET_129),.TB3S(GND),.C3Z(NET_561),.Q3Z(m1_m1_control[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_D12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_432),.B0I1(NET_430),.B0I2(NET_433),.B0I3(NET_431),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T0I0(NET_432),.T0I1(NET_430),.T0I2(NET_433),.T0I3(NET_431),.TB0S(NET_434),.C0Z(NET_422),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_D12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[26]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_control[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D12_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_129),.B2I1(fpgaio_in_int[26]),.B2I2(NET_111),.B2I3(m1_m1_control[26]),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T2I0(NET_129),.T2I1(fpgaio_in_int[22]),.T2I2(NET_111),.T2I3(m1_m1_control[22]),.TB2S(GND),.B2Z(NET_525),.C2Z(NET_433),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_D12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_448),.B3I1(NET_449),.B3I2(NET_451),.B3I3(NET_450),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T3I0(NET_451),.T3I1(NET_450),.T3I2(NET_448),.T3I3(NET_449),.TB3S(NET_452),.C3Z(NET_440),.Q3Z(m1_m1_control[22]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_D14_0 (.tFragBitInfo(16'b0000001100000010),.bFragBitInfo(16'b0000000000000001),.B0I0(apb_fsm[1]),.B0I1(GND),.B0I2(GND),.B0I3(GND),.CD0S(GND),.Q0DI(GND),.Q0EN(nx10146z2),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T0I0(apb_fsm[1]),.T0I1(GND),.T0I2(apb_fsm[0]),.T0I3(lint_WEN_int),.TB0S(GND),.B0Z(not_apb_fsm_1),.Q0Z(apb_fsm[1]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_D14_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(apb_fsm[0]),.T1I2(GND),.T1I3(GND),.TB1S(GND),.C1Z(not_apb_fsm_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_D14_2 (.tFragBitInfo(16'b0011001000010000),.bFragBitInfo(16'b1110111111101110),.B2I0(apb_fsm[1]),.B2I1(apb_fsm[0]),.B2I2(lint_GNT_dup_0),.B2I3(lint_REQ_int),.CD2S(GND),.Q2EN(nx10146z2),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T2I0(apb_fsm[1]),.T2I1(GND),.T2I2(nx10146z1),.T2I3(not_apb_fsm_0),.TB2S(GND),.B2Z(nx10146z2),.Q2Z(apb_fsm[0]),.B2CO(),.C2Z(),.Q2DI(GND),.T2CO());

	LOGIC_3 QL_INST_D14_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_GNT_dup_0),.Q3EN(not_apb_fsm_1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(GND),.T3I2(apb_fsm[0]),.T3I3(lint_WEN_int),.TB3S(GND),.C3Z(nx10146z1),.Q3Z(lint_VALID_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_D15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m1_m1_mode_dup_0[0]),.B0I1(NET_129),.B0I2(NET_128),.B0I3(fpgaio_out_dup_0[76]),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T0I0(m1_m1_mode_dup_0[0]),.T0I1(NET_129),.T0I2(NET_128),.T0I3(fpgaio_out_dup_0[76]),.TB0S(NET_233),.C0Z(NET_230),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_D15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B1I0(m1_m1_control[0]),.B1I1(fpgaio_out_dup_0[64]),.B1I2(NET_128),.B1I3(NET_129),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T1I0(NET_128),.T1I1(NET_129),.T1I2(m1_m1_control[0]),.T1I3(fpgaio_out_dup_0[64]),.TB1S(NET_130),.C1Z(NET_120),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_D15_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0100000000000000),.B2I0(GND),.B2I1(NET_122),.B2I2(NET_120),.B2I3(NET_121),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T2I0(NET_16),.T2I1(lint_ADDR_int[11]),.T2I2(GND),.T2I3(NET_8_CAND5_TLSBL_4_tpGCLKBUF),.TB2S(GND),.B2Z(NET_78),.C2Z(NET_128),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_D15_3 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.T3I0(NET_231),.T3I1(NET_232),.T3I2(GND),.T3I3(NET_230),.TB3S(GND),.C3Z(NET_213),.Q3Z(m1_m1_control[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_D16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx4939z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[44]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[67]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D17_3 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[5]),.T3I1(lint_ADDR_int[3]),.T3I2(lint_ADDR_int[4]),.T3I3(lint_ADDR_int[6]),.C3Z(NET_16),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_D18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[79]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[70]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D18_2 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(NET_30),.T2I2(GND),.T2I3(NET_10),.TB2S(GND),.C2Z(NET_29),.Q2Z(fpgaio_oe_dup_0[68]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_D18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[73]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[76]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[23]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_control[23]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx4939z1_CAND5_BLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[43]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D19_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.T3I0(NET_127),.T3I1(fpgaio_in_int[55]),.T3I2(NET_119),.T3I3(m1_m0_control[23]),.TB3S(GND),.C3Z(NET_452),.Q3Z(fpgaio_oe_dup_0[77]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_D20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[22]),.Q0EN(nx4939z1_CAND5_BLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[54]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx4939z1_CAND5_BLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[47]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[22]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_control[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D22_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.T1I0(NET_119),.T1I1(fpgaio_in_int[54]),.T1I2(NET_127),.T1I3(m1_m0_control[22]),.C1Z(NET_434),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_D22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx9707z1_CAND2_BLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[36]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx4939z1_CAND5_BLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[63]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D23_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[60]),.T2I1(NET_127),.T2I2(NET_119),.T2I3(m1_m0_control[28]),.TB2S(GND),.C2Z(NET_562),.Q2Z(m1_m0_control[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_D23_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_control[26]),.T3I1(NET_127),.T3I2(NET_119),.T3I3(fpgaio_in_int[58]),.TB3S(GND),.C3Z(NET_526),.Q3Z(m1_m0_control[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_D24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx4939z1_CAND5_BLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[38]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_control[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D25_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.T3I0(NET_127),.T3I1(NET_119),.T3I2(fpgaio_in_int[61]),.T3I3(m1_m0_control[29]),.TB3S(GND),.C3Z(NET_580),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_D28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[8]),.Q1EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_waddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[2]),.Q1EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_waddr_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[6]),.Q2EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_waddr_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[11]),.Q3EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_waddr_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[10]),.Q0EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_waddr_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[7]),.Q1EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_waddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[4]),.Q2EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_waddr_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[5]),.Q3EN(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_waddr_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[1]),.Q0EN(nx34006z1_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_waddr_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[0]),.Q1EN(nx34006z1_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_waddr_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[7]),.Q2EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_raddr_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_raddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[5]),.Q0EN(nx34006z1_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_waddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[6]),.Q1EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_raddr_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[5]),.Q2EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_raddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int_11__CAND5_TLSTL_5_tpGCLKBUF),.Q3EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_raddr_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[8]),.Q0EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_raddr_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx44608z1_CAND3_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx44608z1_CAND3_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx44608z1_CAND3_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx44608z1_CAND3_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx39840z1_CAND4_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx39840z1_CAND4_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx39840z1_CAND4_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx39840z1_CAND4_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx39840z1_CAND4_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E11_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_3__CAND3_TLSBL_5_padClk),.QRT(not_RESET_3),.QST(GND),.T0I0(cnt3[0]),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND),.Q0Z(cnt3[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E11_1 (.tFragBitInfo(16'b0000000000010010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_3__CAND3_TLSBL_5_padClk),.QRT(not_RESET_3),.QST(GND),.T1I0(cnt3[0]),.T1I1(GND),.T1I2(cnt3[1]),.T1I3(GND),.TB1S(GND),.Q1Z(cnt3[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E11_2 (.tFragBitInfo(16'b0000000001101100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_3__CAND3_TLSBL_5_padClk),.QRT(not_RESET_3),.QST(GND),.T2I0(cnt3[0]),.T2I1(cnt3[2]),.T2I2(cnt3[1]),.T2I3(GND),.TB2S(GND),.Q2Z(cnt3[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_3__CAND3_TLSBL_5_padClk),.QRT(not_RESET_3),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[22]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.Q0Z(m0_m0_control[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E12_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_in_int[19]),.T1I1(NET_129),.T1I2(m1_m1_control[19]),.T1I3(NET_111),.TB1S(GND),.C1Z(NET_380),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_E12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(cnt3[0]),.B2I1(NET_108),.B2I2(NET_118),.B2I3(m0_m0_control[22]),.CD2S(VCC),.Q2DI(lint_WDATA_int[23]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.T2I0(cnt3[0]),.T2I1(NET_108),.T2I2(NET_118),.T2I3(m0_m0_control[22]),.TB2S(NET_435),.C2Z(NET_431),.Q2Z(m0_m0_control[23]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_E12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B3I0(NET_118),.B3I1(cnt3[1]),.B3I2(m0_m0_control[23]),.B3I3(NET_108),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_control[23]),.T3I1(NET_108),.T3I2(NET_118),.T3I3(cnt3[1]),.TB3S(NET_453),.C3Z(NET_449),.Q3Z(m1_m1_control[19]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_E13_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.T0I0(NET_78),.T0I1(NET_81),.T0I2(NET_80),.T0I3(NET_79),.TB0S(GND),.Q0Z(lint_RDATA_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_524),.B1I1(NET_522),.B1I2(NET_525),.B1I3(NET_523),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.T1I0(NET_525),.T1I1(NET_523),.T1I2(NET_524),.T1I3(NET_522),.TB1S(NET_526),.C1Z(NET_514),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_E13_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.T2I0(NET_213),.T2I1(NET_215),.T2I2(NET_214),.T2I3(NET_216),.TB2S(GND),.Q2Z(lint_RDATA_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E13_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.T3I0(NET_707),.T3I1(NET_705),.T3I2(NET_706),.T3I3(NET_708),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E14_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.T0I0(NET_712),.T0I1(NET_713),.T0I2(NET_711),.T0I3(NET_710),.TB0S(GND),.C0Z(NET_708),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E14_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000001101),.B2I0(apb_fsm[1]),.B2I1(apb_fsm[0]),.B2I2(GND),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.T2I0(nx10146z1),.T2I1(GND),.T2I2(lint_GNT_dup_0),.T2I3(lint_REQ_int),.TB2S(GND),.B2Z(nx7012z3),.C2Z(nx7012z2),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_E14_3 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3EN(nx7012z3),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.T3I0(apb_fsm[1]),.T3I1(apb_fsm[0]),.T3I2(nx7012z2),.T3I3(GND),.TB3S(GND),.Q3Z(lint_GNT_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.Q3DI(GND),.T3CO());

	LOGIC_0 QL_INST_E15_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_221),.B0I1(NET_218),.B0I2(NET_220),.B0I3(NET_219),.T0I0(lint_ADDR_int[16]),.T0I1(lint_ADDR_int[18]),.T0I2(lint_ADDR_int[19]),.T0I3(lint_ADDR_int[17]),.TB0S(GND),.B0Z(NET_216),.C0Z(NET_73),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_E15_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[18]),.T1I1(GND),.T1I2(lint_ADDR_int[19]),.T1I3(lint_ADDR_int[17]),.C1Z(NET_143),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_E15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E15_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_93),.T3I1(NET_92),.T3I2(NET_91),.T3I3(NET_90),.TB3S(GND),.C3Z(NET_81),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_E16_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B0I0(m1_m0_control[7]),.B0I1(NET_119),.B0I2(NET_118),.B0I3(fpgaio_in_int[71]),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.T0I0(NET_97),.T0I1(fpgaio_out_dup_0[44]),.T0I2(i_events[12]),.T0I3(NET_96),.TB0S(GND),.B0Z(NET_466),.C0Z(NET_221),.Q0Z(i_events[0]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(i_events[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E16_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.T2I0(NET_97),.T2I1(fpgaio_out_dup_0[34]),.T2I2(i_events[2]),.T2I3(NET_96),.TB2S(GND),.C2Z(NET_713),.Q2Z(i_events[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_E16_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF),.QST(GND),.T3I0(NET_97),.T3I1(i_events[0]),.T3I2(NET_96),.T3I3(fpgaio_out_dup_0[32]),.TB3S(GND),.C3Z(NET_93),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_E17_0 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T0I0(NET_10),.T0I1(lint_ADDR_int[11]),.T0I2(NET_98),.T0I3(lint_ADDR_int[3]),.TB0S(GND),.C0Z(NET_97),.Q0Z(fpgaio_oe_dup_0[66]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E17_1 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(lint_ADDR_int[5]),.T1I2(lint_ADDR_int[6]),.T1I3(lint_ADDR_int[4]),.C1Z(NET_98),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_E17_2 (.tFragBitInfo(16'b0101111101011111),.bFragBitInfo(16'b0100110001011111),.B2I0(m1_m0_dataout_int[2]),.B2I1(lint_ADDR_int[11]),.B2I2(NET_94_CAND3_BLSTL_5_tpGCLKBUF),.B2I3(fpgaio_oe_dup_0[66]),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T2I0(m1_m0_dataout_int[2]),.T2I1(lint_ADDR_int[11]),.T2I2(NET_94_CAND3_BLSTL_5_tpGCLKBUF),.T2I3(fpgaio_oe_dup_0[66]),.TB2S(NET_20),.C2Z(NET_712),.Q2Z(m0_oper0_wmode_dup_0[1]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_E17_3 (.tFragBitInfo(16'b0000111111111111),.bFragBitInfo(16'b0111011100000111),.B3I0(m1_m0_dataout_int[0]),.B3I1(NET_94_CAND3_BLSTL_5_tpGCLKBUF),.B3I2(fpgaio_oe_dup_0[64]),.B3I3(lint_ADDR_int[11]),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_oe_dup_0[64]),.T3I1(lint_ADDR_int[11]),.T3I2(m1_m0_dataout_int[0]),.T3I3(NET_94_CAND3_BLSTL_5_tpGCLKBUF),.TB3S(NET_20),.C3Z(NET_92),.Q3Z(m1_m0_control[7]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_E18_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_oe_dup_0[73]),.B0I1(NET_21),.B0I2(NET_20),.B0I3(i_events[9]),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T0I0(NET_127),.T0I1(m1_m0_control[21]),.T0I2(fpgaio_in_int[53]),.T0I3(NET_119),.TB0S(GND),.B0Z(NET_152),.C0Z(NET_416),.Q0Z(m1_m0_control[21]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[9]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(i_events[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[72]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[72]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E19_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T0I0(NET_20),.T0I1(fpgaio_oe_dup_0[69]),.T0I2(i_events[5]),.T0I3(NET_21),.TB0S(GND),.C0Z(NET_647),.Q0Z(fpgaio_oe_dup_0[75]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E19_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(NET_21),.T1I1(NET_20),.T1I2(i_events[14]),.T1I3(fpgaio_oe_dup_0[78]),.TB1S(GND),.C1Z(NET_254),.Q1Z(i_events[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_E19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E19_3 (.tFragBitInfo(16'b0101010111111111),.bFragBitInfo(16'b0010101000111111),.B3I0(lint_ADDR_int[11]),.B3I1(NET_94_CAND3_BLSTL_5_tpGCLKBUF),.B3I2(m1_m0_dataout_int[12]),.B3I3(fpgaio_oe_dup_0[76]),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_dataout_int[12]),.T3I1(fpgaio_oe_dup_0[76]),.T3I2(lint_ADDR_int[11]),.T3I3(NET_94_CAND3_BLSTL_5_tpGCLKBUF),.TB3S(NET_20),.C3Z(NET_220),.Q3Z(i_events[5]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_E20_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx4939z1_CAND5_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T0I0(m1_m0_control[24]),.T0I1(NET_119),.T0I2(NET_127),.T0I3(fpgaio_in_int[56]),.TB0S(GND),.C0Z(NET_491),.Q0Z(fpgaio_out_dup_0[62]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx4939z1_CAND5_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[34]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_control[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx4939z1_CAND5_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[57]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx4939z1_CAND5_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[32]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx4939z1_CAND5_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[37]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx4939z1_CAND5_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[39]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx4939z1_CAND5_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[59]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_control[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E24_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T2I0(NET_119),.T2I1(fpgaio_in_int[51]),.T2I2(m1_m0_control[19]),.T2I3(NET_127),.TB2S(GND),.C2Z(NET_381),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_E24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx9707z1_CAND2_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[45]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E25_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.T0I0(NET_119),.T0I1(m1_m0_clr_dup_0),.T0I2(fpgaio_in_int[49]),.T0I3(NET_127),.TB0S(GND),.C0Z(NET_344),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_E25_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_119),.T1I1(fpgaio_in_int[50]),.T1I2(m1_m0_sat_dup_0),.T1I3(NET_127),.TB1S(GND),.C1Z(NET_362),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_E25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx9707z1_CAND2_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[47]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(m1_m0_clr_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx22245z1_CAND3_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[8]),.Q2EN(nx60831z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_raddr_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[11]),.Q0EN(nx60831z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_raddr_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[6]),.Q1EN(nx60831z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_raddr_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[3]),.Q2EN(nx60831z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_raddr_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx22245z1_CAND3_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[1]),.Q0EN(nx22245z1_CAND3_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_waddr_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[4]),.Q1EN(nx60831z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_raddr_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[9]),.Q2EN(nx60831z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_raddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx60831z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_raddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[9]),.Q0EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_raddr_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[1]),.Q1EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_raddr_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[3]),.Q2EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_raddr_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[0]),.Q3EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_raddr_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(NET_762),.Q0EN(nx34006z1_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_we_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[2]),.Q1EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_raddr_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[4]),.Q3EN(nx34850z1),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_raddr_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx44608z1_CAND3_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000010000000),.B2I0(lint_ADDR_int[12]),.B2I1(NET_144),.B2I2(NET_65),.B2I3(lint_ADDR_int[13]),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B2Z(nx34006z1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx44608z1_CAND3_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx39840z1_CAND4_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F6_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0001000000000000),.B2I0(lint_ADDR_int[13]),.B2I1(lint_ADDR_int[14]),.B2I2(lint_ADDR_int[12]),.B2I3(lint_WEN_int),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(NET_367),.T2I1(NET_142),.T2I2(NET_141),.T2I3(GND),.TB2S(GND),.B2Z(NET_367),.C2Z(nx34850z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_F6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx39840z1_CAND4_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F7_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx39840z1_CAND4_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(NET_60),.T2I1(m0_oper0_wmode_dup_0[1]),.T2I2(fpgaio_out_dup_0[3]),.T2I3(NET_61),.TB2S(GND),.C2Z(NET_703),.Q2Z(fpgaio_out_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_F7_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx39840z1_CAND4_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(NET_60),.T3I1(fpgaio_out_dup_0[1]),.T3I2(m0_oper0_rmode_dup_0[1]),.T3I3(NET_61),.TB3S(GND),.C3Z(NET_56),.Q3Z(fpgaio_out_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_F8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000010000000000),.B0I0(GND),.B0I1(NET_8),.B0I2(GND),.B0I3(NET_30),.B0Z(NET_58),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m0_m0_clr_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F10_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_102),.B0I1(fpgaio_out_dup_0[19]),.B0I2(m1_ram_control[19]),.B0I3(NET_85),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_out_dup_0[15]),.T0I1(NET_61),.T0I2(m0_ram_control[15]),.T0I3(NET_60),.TB0S(GND),.B0Z(NET_375),.C0Z(NET_309),.Q0Z(m1_ram_control[21]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(m0_ram_control[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_102),.B2I1(fpgaio_out_dup_0[21]),.B2I2(NET_85),.B2I3(m1_ram_control[21]),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.B2Z(NET_410),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F10_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(NET_67),.T3I1(NET_65),.T3I2(NET_68),.T3I3(lint_ADDR_int[6]),.C3Z(nx44608z1),.Q3Z(m1_ram_control[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_F11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_576),.B1I1(NET_578),.B1I2(NET_579),.B1I3(NET_577),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T1I0(NET_579),.T1I1(NET_577),.T1I2(NET_576),.T1I3(NET_578),.TB1S(NET_580),.C1Z(NET_568),.Q1Z(m1_ram_control[24]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_F11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F11_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_out_dup_0[24]),.T3I1(NET_85),.T3I2(m1_ram_control[24]),.T3I3(NET_102),.C3Z(NET_485),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_F12_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.T0I0(NET_459),.T0I1(NET_460),.T0I2(NET_457),.T0I3(NET_458),.TB0S(GND),.Q0Z(lint_RDATA_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_559),.B1I1(NET_560),.B1I2(NET_558),.B1I3(NET_561),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.T1I0(NET_558),.T1I1(NET_561),.T1I2(NET_559),.T1I3(NET_560),.TB1S(NET_562),.C1Z(NET_550),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_F12_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.T2I0(m1_m1_sat_dup_0),.T2I1(NET_111),.T2I2(NET_129),.T2I3(fpgaio_in_int[18]),.TB2S(GND),.C2Z(NET_361),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_F12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_361),.B3I1(NET_359),.B3I2(NET_358),.B3I3(NET_360),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.T3I0(NET_358),.T3I1(NET_360),.T3I2(NET_361),.T3I3(NET_359),.TB3S(NET_362),.C3Z(NET_350),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_F13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(cnt3[2]),.B0I1(NET_108),.B0I2(m0_m0_control[24]),.B0I3(NET_118),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T0I0(cnt3[2]),.T0I1(NET_108),.T0I2(m0_m0_control[24]),.T0I3(NET_118),.TB0S(NET_492),.C0Z(NET_488),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_490),.B1I1(NET_487),.B1I2(NET_488),.B1I3(NET_489),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T1I0(NET_488),.T1I1(NET_489),.T1I2(NET_490),.T1I3(NET_487),.TB1S(NET_491),.C1Z(NET_479),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_F13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m0_m0_control[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_379),.B3I1(NET_377),.B3I2(NET_378),.B3I3(NET_380),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(NET_378),.T3I1(NET_380),.T3I2(NET_379),.T3I3(NET_377),.TB3S(NET_381),.C3Z(NET_369),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_F14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000100),.B0I0(lint_GNT_dup_0),.B0I1(lint_REQ_int),.B0I2(apb_fsm[0]),.B0I3(apb_fsm[1]),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(GND),.B0Z(NET_142),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F14_1 (.tFragBitInfo(16'b0000000000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_REQ_int),.Q1EN(RESET_int[0]),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(GND),.T1I0(apb_fsm[0]),.T1I1(GND),.T1I2(GND),.T1I3(apb_fsm[1]),.TB1S(GND),.C1Z(NET_65),.Q1Z(saved_REQ),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_F14_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_464),.B2I1(NET_463),.B2I2(NET_465),.B2I3(NET_462),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(GND),.T2I0(NET_37),.T2I1(NET_60),.T2I2(fpgaio_out_dup_0[31]),.T2I3(saved_REQ),.TB2S(GND),.B2Z(NET_460),.C2Z(NET_616),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_F14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F15_0 (.tFragBitInfo(16'b0010000000100011),.bFragBitInfo(16'b0000000000000010),.B0I0(NET_143),.B0I1(lint_ADDR_int[15]),.B0I2(lint_ADDR_int[16]),.B0I3(lint_ADDR_int[14]),.T0I0(lint_ADDR_int[14]),.T0I1(GND),.T0I2(lint_ADDR_int[13]),.T0I3(lint_ADDR_int[12]),.TB0S(GND),.B0Z(NET_144),.C0Z(NET_620),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_F15_1 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[14]),.T1I1(lint_ADDR_int[15]),.T1I2(lint_ADDR_int[16]),.T1I3(lint_ADDR_int[12]),.C1Z(NET_253),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_F15_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000000000010),.B2I0(NET_143),.B2I1(lint_ADDR_int[15]),.B2I2(lint_ADDR_int[16]),.B2I3(GND),.T2I0(NET_142),.T2I1(lint_WEN_int),.T2I2(NET_171),.T2I3(lint_ADDR_int[13]),.TB2S(GND),.B2Z(NET_141),.C2Z(nx60831z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_F15_3 (.tFragBitInfo(16'b1100000000000000),.bFragBitInfo(16'b1000110000000000),.B3I0(NET_171),.B3I1(apb_fsm[1]),.B3I2(NET_620),.B3I3(apb_fsm[0]),.T3I0(NET_620),.T3I1(apb_fsm[0]),.T3I2(NET_171),.T3I3(apb_fsm[1]),.TB3S(NET_141),.C3Z(NET_621),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_F16_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_out_dup_0[39]),.T0I1(NET_97),.T0I2(i_events[7]),.T0I3(NET_96),.TB0S(GND),.C0Z(NET_465),.Q0Z(i_events[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F16_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T1I0(i_events[6]),.T1I1(NET_97),.T1I2(fpgaio_out_dup_0[38]),.T1I3(NET_96),.TB1S(GND),.C1Z(NET_631),.Q1Z(m0_m0_outsel_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_F16_2 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_118),.B2I1(fpgaio_in_int[64]),.B2I2(m1_m0_outsel_dup_0[0]),.B2I3(NET_119),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T2I0(NET_67),.T2I1(NET_602),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(NET_104),.C2Z(nx9707z1),.Q2Z(i_events[7]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_F16_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_in_int[66]),.T3I1(NET_119),.T3I2(m1_m0_outsel_dup_0[2]),.T3I3(NET_118),.C3Z(NET_714),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_F17_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000001000000000),.B0I0(NET_22),.B0I1(GND),.B0I2(GND),.B0I3(NET_8),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T0I0(i_events[3]),.T0I1(NET_20),.T0I2(NET_21),.T0I3(fpgaio_oe_dup_0[67]),.TB0S(GND),.B0Z(NET_37),.C0Z(NET_686),.Q0Z(i_events[3]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_65),.B1I1(lint_ADDR_int[3]),.B1I2(NET_68),.B1I3(lint_ADDR_int[4]),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(NET_68),.T1I1(lint_ADDR_int[4]),.T1I2(NET_65),.T1I3(lint_ADDR_int[3]),.TB1S(lint_ADDR_int[6]),.C1Z(nx58292z1),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_F17_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0100000000000000),.B2I0(lint_ADDR_int[4]),.B2I1(lint_ADDR_int[6]),.B2I2(lint_ADDR_int[5]),.B2I3(lint_ADDR_int[3]),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(NET_22),.T2I1(GND),.T2I2(lint_ADDR_int[11]),.T2I3(NET_8),.TB2S(GND),.B2Z(NET_22),.C2Z(NET_118),.Q2Z(fpgaio_out_dup_0[65]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_F17_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(NET_10),.T3I1(NET_22),.T3I2(GND),.T3I3(GND),.TB3S(GND),.C3Z(NET_21),.Q3Z(fpgaio_oe_dup_0[65]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_F18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_20),.B0I1(NET_21),.B0I2(i_events[1]),.B0I3(fpgaio_oe_dup_0[65]),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0Z(NET_0),.Q0Z(i_events[4]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F18_1 (.tFragBitInfo(16'b0101010111111111),.bFragBitInfo(16'b0011111100010101),.B1I0(fpgaio_oe_dup_0[71]),.B1I1(NET_94_CAND3_BLSTL_6_tpGCLKBUF),.B1I2(m1_m0_dataout_int[7]),.B1I3(lint_ADDR_int[11]),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(m1_m0_dataout_int[7]),.T1I1(lint_ADDR_int[11]),.T1I2(fpgaio_oe_dup_0[71]),.T1I3(NET_94_CAND3_BLSTL_6_tpGCLKBUF),.TB1S(NET_20),.C1Z(NET_464),.Q1Z(fpgaio_out_dup_0[78]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_F18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q2Z(i_events[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F18_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_oe_dup_0[68]),.T3I1(NET_20),.T3I2(NET_21),.T3I3(i_events[4]),.TB3S(GND),.C3Z(NET_667),.Q3Z(fpgaio_oe_dup_0[74]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_F19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(i_events[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F19_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_oe_dup_0[75]),.T1I1(NET_21),.T1I2(i_events[11]),.T1I3(NET_20),.TB1S(GND),.C1Z(NET_194),.Q1Z(i_events[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_F19_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(NET_20),.T2I1(NET_21),.T2I2(fpgaio_oe_dup_0[77]),.T2I3(i_events[13]),.TB2S(GND),.C2Z(NET_234),.Q2Z(fpgaio_oe_dup_0[79]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_F19_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(NET_20),.T3I1(NET_21),.T3I2(fpgaio_oe_dup_0[79]),.T3I3(i_events[15]),.C3Z(NET_292),.Q3Z(i_events[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_F20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(m1_m1_tc_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx4939z1_CAND5_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[41]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx4939z1_CAND5_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[51]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_outsel_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx4939z1_CAND5_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[45]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx4939z1_CAND5_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[35]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[8]),.Q1EN(nx9707z1_CAND2_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[40]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx9707z1_CAND2_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[33]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_outsel_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx9707z1_CAND2_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[43]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F27_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_65),.T1I1(lint_ADDR_int[13]),.T1I2(NET_171),.T1I3(GND),.C1Z(nx22245z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_F27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[18]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_sat_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(NET_762),.Q0EN(nx22245z1_CAND3_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_we_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[3]),.Q1EN(nx22245z1_CAND3_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_waddr_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[2]),.Q2EN(nx60831z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_raddr_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F31_3 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1110000011101111),.B3I0(lint_ADDR_int[13]),.B3I1(lint_ADDR_int[12]),.B3I2(apb_fsm[0]),.B3I3(lint_ADDR_int[11]),.CD3S(VCC),.Q3DI(lint_ADDR_int[0]),.Q3EN(nx22245z1_CAND3_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(apb_fsm[0]),.T3I1(lint_ADDR_int[11]),.T3I2(lint_ADDR_int[13]),.T3I3(lint_ADDR_int[12]),.TB3S(m1_oper0_rdata_int[30]),.C3Z(NET_750),.Q3Z(m1_oper0_waddr_dup_0[0]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_F32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[5]),.Q0EN(nx60831z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_raddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[0]),.Q1EN(nx60831z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_raddr_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[1]),.Q2EN(nx60831z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_raddr_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[7]),.Q3EN(nx60831z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_raddr_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(m0_m0_dataout_int[1]),.B0I1(NET_58),.B0I2(NET_59),.B0I3(fpgaio_oe_dup_0[1]),.B0Z(NET_55),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G5_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(fpgaio_oe_dup_0[15]),.T3I1(m0_m0_dataout_int[15]),.T3I2(NET_58),.T3I3(NET_59),.C3Z(NET_308),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx39840z1_CAND4_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx39840z1_CAND4_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G7_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_56),.T2I1(NET_54),.T2I2(NET_55),.T2I3(NET_53),.TB2S(GND),.C2Z(NET_57),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_G7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx39840z1_CAND4_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.Q2Z(m0_m0_osel_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G8_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.T3I0(apb_fsm[0]),.T3I1(lint_ADDR_int[2]),.T3I2(lint_ADDR_int[7]),.T3I3(lint_ADDR_int[8]),.C3Z(NET_8),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[29]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[18]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.Q2Z(m0_m0_sat_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G10_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T0I0(NET_309),.T0I1(NET_306),.T0I2(NET_308),.T0I3(NET_307),.TB0S(GND),.C0Z(NET_310),.Q0Z(m1_ram_control[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G10_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[6]),.T1I1(NET_146),.T1I2(NET_68),.T1I3(NET_65),.C1Z(nx39840z1),.Q1Z(m1_ram_control[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_102),.B2I1(NET_85),.B2I2(fpgaio_out_dup_0[26]),.B2I3(m1_ram_control[26]),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.B2Z(NET_520),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G10_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(NET_102),.T3I1(NET_85),.T3I2(m1_ram_control[28]),.T3I3(fpgaio_out_dup_0[28]),.TB3S(GND),.C3Z(NET_556),.Q3Z(m0_oper1_wmode_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_G11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.Q0Z(m1_ram_control[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G11_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(NET_102),.T1I1(NET_85),.T1I2(m1_ram_control[29]),.T1I3(fpgaio_out_dup_0[29]),.C1Z(NET_574),.Q1Z(m1_ram_control[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_85),.B2I1(fpgaio_out_dup_0[17]),.B2I2(m1_ram_control[17]),.B2I3(NET_102),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.B2Z(NET_338),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G11_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(NET_102),.T3I1(NET_85),.T3I2(fpgaio_out_dup_0[18]),.T3I3(m1_ram_control[18]),.C3Z(NET_356),.Q3Z(m1_ram_control[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G12_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.T0I0(NET_552),.T0I1(NET_551),.T0I2(NET_550),.T0I3(NET_549),.TB0S(GND),.Q0Z(lint_RDATA_dup_0[28]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_341),.B1I1(NET_343),.B1I2(NET_340),.B1I3(NET_342),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.T1I0(NET_340),.T1I1(NET_342),.T1I2(NET_341),.T1I3(NET_343),.TB1S(NET_344),.C1Z(NET_331),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_G12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m0_m0_clr_dup_0),.B2I1(NET_108),.B2I2(cnt1[1]),.B2I3(NET_118),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.T2I0(m0_m0_clr_dup_0),.T2I1(NET_108),.T2I2(cnt1[1]),.T2I3(NET_118),.TB2S(NET_345),.C2Z(NET_341),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_G12_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.T3I0(m1_m1_clr_dup_0),.T3I1(NET_129),.T3I2(fpgaio_in_int[17]),.T3I3(NET_111),.TB3S(GND),.C3Z(NET_343),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_G13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_415),.B0I1(NET_414),.B0I2(NET_412),.B0I3(NET_413),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.T0I0(NET_415),.T0I1(NET_414),.T0I2(NET_412),.T0I3(NET_413),.TB0S(NET_416),.C0Z(NET_404),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G13_1 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.T1I0(NET_624),.T1I1(NET_626),.T1I2(NET_623),.T1I3(NET_625),.TB1S(GND),.Q1Z(lint_RDATA_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_G13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_520),.B2I1(NET_518),.B2I2(GND),.B2I3(NET_519),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.B2Z(NET_516),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G13_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.T3I0(NET_515),.T3I1(NET_513),.T3I2(NET_516),.T3I3(NET_514),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_G14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m0_m0_control[26]),.B0I1(NET_108),.B0I2(NET_118),.B0I3(cnt4[1]),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T0I0(m0_m0_control[26]),.T0I1(NET_108),.T0I2(NET_118),.T0I3(cnt4[1]),.TB0S(NET_527),.C0Z(NET_523),.Q0Z(m0_m0_control[26]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G14_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(m0_oper1_wmode_dup_0[1]),.T1I1(fpgaio_out_dup_0[7]),.T1I2(NET_102),.T1I3(NET_103),.TB1S(GND),.C1Z(NET_462),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_G14_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_409),.B2I1(NET_410),.B2I2(GND),.B2I3(NET_408),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T2I0(m0_oper1_wmode_dup_0[0]),.T2I1(fpgaio_out_dup_0[6]),.T2I2(NET_102),.T2I3(NET_103),.TB2S(GND),.B2Z(NET_406),.C2Z(NET_628),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_G14_3 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_555),.T3I2(NET_554),.T3I3(NET_556),.C3Z(NET_552),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G15_0 (.tFragBitInfo(16'b0001010001000100),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_60),.B0I1(cnt4[2]),.B0I2(fpgaio_out_dup_0[27]),.B0I3(NET_37),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_4__CAND4_TLSBL_7_padClk),.QRT(not_RESET_1),.QST(GND),.T0I0(GND),.T0I1(cnt4[2]),.T0I2(cnt4[0]),.T0I3(cnt4[1]),.TB0S(GND),.B0Z(NET_545),.Q0Z(cnt4[2]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G15_1 (.tFragBitInfo(16'b0000000100010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_4__CAND4_TLSBL_7_padClk),.QRT(not_RESET_1),.QST(GND),.T1I0(GND),.T1I1(GND),.T1I2(cnt4[0]),.T1I3(cnt4[1]),.TB1S(GND),.Q1Z(cnt4[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_G15_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000001000000000),.B2I0(NET_31),.B2I1(lint_ADDR_int[11]),.B2I2(GND),.B2I3(NET_10),.QCK(CLK_int_4__CAND4_TLSBL_7_padClk),.QRT(not_RESET_1),.QST(GND),.T2I0(NET_628),.T2I1(NET_631),.T2I2(NET_629),.T2I3(NET_630),.TB2S(GND),.B2Z(NET_129),.C2Z(NET_626),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_G15_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_4__CAND4_TLSBL_7_padClk),.QRT(not_RESET_1),.QST(GND),.T3I0(GND),.T3I1(GND),.T3I2(cnt4[0]),.T3I3(GND),.TB3S(GND),.Q3Z(cnt4[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_G16_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T0I0(NET_36),.T0I1(NET_37),.T0I2(fpgaio_in_int[65]),.T0I3(m0_m0_outsel_dup_0[1]),.TB0S(GND),.C0Z(NET_23),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G16_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(NET_36),.T1I1(NET_37),.T1I2(m0_m0_outsel_dup_0[3]),.T1I3(fpgaio_in_int[67]),.TB1S(GND),.C1Z(NET_691),.Q1Z(m0_m0_control[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_G16_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B2I0(fpgaio_in_int[75]),.B2I1(NET_37),.B2I2(NET_36),.B2I3(m0_m0_control[11]),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T2I0(NET_118),.T2I1(fpgaio_in_int[70]),.T2I2(NET_119),.T2I3(m1_m0_tc_dup_0),.TB2S(GND),.B2Z(NET_199),.C2Z(NET_632),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_G16_3 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(lint_ADDR_int[11]),.T3I2(NET_8_CAND5_TLSBL_7_tpGCLKBUF),.T3I3(NET_31),.C3Z(NET_119),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G17_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000001000000000),.B0I0(NET_16),.B0I1(GND),.B0I2(GND),.B0I3(NET_8),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[3]),.T0I1(lint_ADDR_int[4]),.T0I2(NET_9),.T0I3(NET_8),.TB0S(GND),.B0Z(NET_12),.C0Z(NET_20),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G17_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(NET_118),.T1I1(m1_m0_mode_dup_0[0]),.T1I2(NET_119),.T1I3(fpgaio_in_int[76]),.C1Z(NET_222),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G17_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(NET_103),.T2I1(m1_m0_dataout_int[21]),.T2I2(m0_ram_control[21]),.T2I3(NET_94_CAND3_BLSTL_7_tpGCLKBUF),.TB2S(GND),.C2Z(NET_409),.Q2Z(m0_ram_control[21]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_G17_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_in_int[78]),.T3I1(NET_37),.T3I2(NET_36),.T3I3(m0_m0_osel_dup_0),.TB3S(GND),.C3Z(NET_259),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_G18_0 (.tFragBitInfo(16'b0111011101110111),.bFragBitInfo(16'b0111000001110111),.B0I0(NET_94_CAND3_BLSTL_7_tpGCLKBUF),.B0I1(m1_m0_dataout_int[6]),.B0I2(lint_ADDR_int[11]),.B0I3(fpgaio_oe_dup_0[70]),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T0I0(NET_94_CAND3_BLSTL_7_tpGCLKBUF),.T0I1(m1_m0_dataout_int[6]),.T0I2(lint_ADDR_int[11]),.T0I3(fpgaio_oe_dup_0[70]),.TB0S(NET_20),.C0Z(NET_630),.Q0Z(i_events[8]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G18_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_oe_dup_0[72]),.T1I1(NET_20),.T1I2(NET_21),.T1I3(i_events[8]),.C1Z(NET_273),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G18_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000010000000000),.B2I0(GND),.B2I1(NET_10),.B2I2(GND),.B2I3(NET_31),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(i_events[10]),.T2I1(NET_20),.T2I2(NET_21),.T2I3(fpgaio_oe_dup_0[74]),.TB2S(GND),.B2Z(NET_28),.C2Z(NET_175),.Q2Z(i_events[10]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_G18_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_dataout_int[30]),.T3I1(NET_5),.T3I2(fpgaio_out_dup_0[62]),.T3I3(NET_59),.TB3S(GND),.C3Z(NET_590),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_G19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(m0_m0_dataout_int[31]),.B0I1(fpgaio_out_dup_0[63]),.B0I2(NET_5),.B0I3(NET_59),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B0Z(NET_608),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G19_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_29_CAND4_BLSTL_7_tpGCLKBUF),.B2I1(fpgaio_oe_dup_0[40]),.B2I2(m1_m1_control[8]),.B2I3(NET_28),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(m0_ram_control[28]),.T2I1(NET_94_CAND3_BLSTL_7_tpGCLKBUF),.T2I2(m1_m0_dataout_int[28]),.T2I3(NET_103),.TB2S(GND),.B2Z(NET_280),.C2Z(NET_555),.Q2Z(m0_ram_control[28]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_G19_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_dataout_int[27]),.T3I1(fpgaio_out_dup_0[59]),.T3I2(NET_5),.T3I3(NET_59),.TB3S(GND),.C3Z(NET_537),.Q3Z(m1_m1_control[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_G20_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_oe_dup_0[43]),.T0I1(NET_28),.T0I2(NET_29_CAND4_BLSTL_7_tpGCLKBUF),.T0I3(m1_m1_control[11]),.TB0S(GND),.C0Z(NET_201),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G20_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_oe_dup_0[36]),.T1I1(NET_28),.T1I2(m1_m1_control[4]),.T1I3(NET_29_CAND4_BLSTL_7_tpGCLKBUF),.TB1S(GND),.C1Z(NET_674),.Q1Z(m1_m1_control[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_G20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_control[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx4939z1_CAND5_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[50]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G21_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T3I0(NET_103),.T3I1(m1_m0_dataout_int[26]),.T3I2(m0_ram_control[26]),.T3I3(NET_94_CAND3_BLSTL_7_tpGCLKBUF),.TB3S(GND),.C3Z(NET_519),.Q3Z(m0_ram_control[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_G22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(m1_m1_control[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G22_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_control[5]),.T1I1(NET_29_CAND4_BLSTL_7_tpGCLKBUF),.T1I2(fpgaio_oe_dup_0[37]),.T1I3(NET_28),.TB1S(GND),.C1Z(NET_654),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_G22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[20]),.Q2EN(nx4939z1_CAND5_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[52]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx4939z1_CAND5_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[60]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx4939z1_CAND5_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[49]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx4939z1_CAND5_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[40]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_osel_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G31_1 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1110000011101111),.B1I0(lint_ADDR_int[13]),.B1I1(lint_ADDR_int[12]),.B1I2(apb_fsm[0]),.B1I3(lint_ADDR_int[11]),.T1I0(apb_fsm[0]),.T1I1(lint_ADDR_int[11]),.T1I2(lint_ADDR_int[13]),.T1I3(lint_ADDR_int[12]),.TB1S(m1_oper0_rdata_int[27]),.C1Z(NET_748),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_G31_2 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1011101110110001),.B2I0(apb_fsm[0]),.B2I1(lint_ADDR_int[11]),.B2I2(lint_ADDR_int[13]),.B2I3(lint_ADDR_int[12]),.T2I0(apb_fsm[0]),.T2I1(lint_ADDR_int[11]),.T2I2(lint_ADDR_int[13]),.T2I3(lint_ADDR_int[12]),.TB2S(m1_oper0_rdata_int[20]),.C2Z(NET_744),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_G31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H2_0 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1011101110110001),.B0I0(apb_fsm[0]),.B0I1(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.B0I2(lint_ADDR_int[13]),.B0I3(lint_ADDR_int[14]),.T0I0(apb_fsm[0]),.T0I1(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.T0I2(lint_ADDR_int[13]),.T0I3(lint_ADDR_int[14]),.TB0S(m0_oper0_rdata_int[15]),.C0Z(NET_305),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_H2_1 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1110000011101111),.B1I0(lint_ADDR_int[13]),.B1I1(lint_ADDR_int[14]),.B1I2(apb_fsm[0]),.B1I3(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.T1I0(apb_fsm[0]),.T1I1(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.T1I2(lint_ADDR_int[13]),.T1I3(lint_ADDR_int[14]),.TB1S(m0_oper0_rdata_int[8]),.C1Z(NET_286),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_H2_2 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1101110111010001),.B2I0(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.B2I1(apb_fsm[0]),.B2I2(lint_ADDR_int[13]),.B2I3(lint_ADDR_int[14]),.T2I0(apb_fsm[0]),.T2I1(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.T2I2(lint_ADDR_int[13]),.T2I3(lint_ADDR_int[14]),.TB2S(m0_oper0_rdata_int[9]),.C2Z(NET_165),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_H2_3 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1110000011101111),.B3I0(lint_ADDR_int[13]),.B3I1(lint_ADDR_int[14]),.B3I2(apb_fsm[0]),.B3I3(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.T3I0(apb_fsm[0]),.T3I1(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.T3I2(lint_ADDR_int[13]),.T3I3(lint_ADDR_int[14]),.TB3S(m0_oper0_rdata_int[10]),.C3Z(NET_188),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_H3_0 (.tFragBitInfo(16'b1010101011111111),.bFragBitInfo(16'b1010100011111101),.B0I0(apb_fsm[0]),.B0I1(lint_ADDR_int[14]),.B0I2(lint_ADDR_int[13]),.B0I3(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.T0I0(apb_fsm[0]),.T0I1(lint_ADDR_int[14]),.T0I2(lint_ADDR_int[13]),.T0I3(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.TB0S(m0_oper0_rdata_int[11]),.C0Z(NET_207),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_H3_1 (.tFragBitInfo(16'b1010101011111111),.bFragBitInfo(16'b1111001110100011),.B1I0(lint_ADDR_int[13]),.B1I1(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.B1I2(apb_fsm[0]),.B1I3(lint_ADDR_int[14]),.T1I0(apb_fsm[0]),.T1I1(lint_ADDR_int[14]),.T1I2(lint_ADDR_int[13]),.T1I3(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.TB1S(m0_oper0_rdata_int[13]),.C1Z(NET_247),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_H3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H3_3 (.tFragBitInfo(16'b1010101011111111),.bFragBitInfo(16'b1111001110100011),.B3I0(lint_ADDR_int[13]),.B3I1(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.B3I2(apb_fsm[0]),.B3I3(lint_ADDR_int[14]),.T3I0(apb_fsm[0]),.T3I1(lint_ADDR_int[14]),.T3I2(lint_ADDR_int[13]),.T3I3(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.TB3S(m0_oper0_rdata_int[14]),.C3Z(NET_267),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_H4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H4_1 (.tFragBitInfo(16'b1111000011111111),.bFragBitInfo(16'b1011101110110001),.B1I0(apb_fsm[0]),.B1I1(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.B1I2(lint_ADDR_int[14]),.B1I3(lint_ADDR_int[13]),.T1I0(lint_ADDR_int[14]),.T1I1(lint_ADDR_int[13]),.T1I2(apb_fsm[0]),.T1I3(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF),.TB1S(m0_oper0_rdata_int[1]),.C1Z(NET_47),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_H4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H10_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.QST(GND),.T0I0(NET_85),.T0I1(fpgaio_out_dup_0[22]),.T0I2(m1_ram_control[22]),.T0I3(NET_102),.TB0S(GND),.C0Z(NET_428),.Q0Z(m0_m0_outsel_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[23]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.QST(GND),.Q2Z(m1_ram_control[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H10_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.QST(GND),.T3I0(NET_85),.T3I1(fpgaio_out_dup_0[23]),.T3I2(m1_ram_control[23]),.T3I3(NET_102),.C3Z(NET_446),.Q3Z(m1_ram_control[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H11_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0100000000000000),.B0I0(GND),.B0I1(NET_445),.B0I2(NET_446),.B0I3(NET_444),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.T0I0(NET_441),.T0I1(NET_442),.T0I2(NET_440),.T0I3(NET_439),.TB0S(GND),.B0Z(NET_442),.Q0Z(lint_RDATA_dup_0[23]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H11_1 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.T1I0(NET_569),.T1I1(NET_567),.T1I2(NET_568),.T1I3(NET_570),.TB1S(GND),.Q1Z(lint_RDATA_dup_0[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H11_3 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.T3I0(GND),.T3I1(NET_572),.T3I2(NET_574),.T3I3(NET_573),.C3Z(NET_570),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H12_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.T0I0(NET_421),.T0I1(NET_422),.T0I2(NET_424),.T0I3(NET_423),.TB0S(GND),.Q0Z(lint_RDATA_dup_0[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B1I0(NET_108),.B1I1(cnt1[2]),.B1I2(NET_118),.B1I3(m0_m0_sat_dup_0),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.T1I0(NET_118),.T1I1(m0_m0_sat_dup_0),.T1I2(NET_108),.T1I3(cnt1[2]),.TB1S(NET_363),.C1Z(NET_359),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_H12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_88),.B2I1(lint_ADDR_int[5]),.B2I2(lint_ADDR_int[6]),.B2I3(NET_10),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.B2Z(NET_85),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H12_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_727),.B3I1(NET_27),.B3I2(NET_42),.B3I3(NET_4),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.T3I0(NET_42),.T3I1(NET_4),.T3I2(NET_727),.T3I3(NET_27),.TB3S(NET_57),.Q3Z(lint_RDATA_dup_0[1]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_H13_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0100000000000000),.B0I0(GND),.B0I1(NET_483),.B0I2(NET_484),.B0I3(NET_485),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.T0I0(NET_404),.T0I1(NET_403),.T0I2(NET_405),.T0I3(NET_406),.TB0S(GND),.B0Z(NET_481),.Q0Z(lint_RDATA_dup_0[21]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H13_1 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.T1I0(NET_369),.T1I1(NET_368),.T1I2(NET_370),.T1I3(NET_371),.TB1S(GND),.Q1Z(lint_RDATA_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H13_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.T2I0(NET_426),.T2I1(NET_427),.T2I2(GND),.T2I3(NET_428),.TB2S(GND),.C2Z(NET_424),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_H13_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.T3I0(NET_478),.T3I1(NET_481),.T3I2(NET_479),.T3I3(NET_480),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_H14_0 (.tFragBitInfo(16'b0000000001101100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T0I0(cnt1[0]),.T0I1(cnt1[2]),.T0I2(cnt1[1]),.T0I3(GND),.TB0S(GND),.Q0Z(cnt1[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H14_1 (.tFragBitInfo(16'b0000000000010010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T1I0(cnt1[0]),.T1I1(GND),.T1I2(cnt1[1]),.T1I3(GND),.TB1S(GND),.Q1Z(cnt1[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H14_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0010000000000000),.B2I0(NET_8_CAND5_TLSBL_8_tpGCLKBUF),.B2I1(GND),.B2I2(NET_88),.B2I3(NET_9),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T2I0(cnt1[0]),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(NET_102),.Q2Z(cnt1[0]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_H14_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T3I0(NET_37),.T3I1(NET_60),.T3I2(cnt1[0]),.T3I3(fpgaio_out_dup_0[16]),.C3Z(NET_326),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H15_0 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000000000000),.T0I0(NET_10),.T0I1(NET_88),.T0I2(NET_9),.T0I3(GND),.TB0S(GND),.C0Z(NET_96),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_H15_1 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(GND),.T1I1(NET_374),.T1I2(NET_375),.T1I3(NET_373),.C1Z(NET_371),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_H15_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0010000000000000),.B2I0(NET_8_CAND5_TLSBL_8_tpGCLKBUF),.B2I1(lint_ADDR_int[6]),.B2I2(NET_88),.B2I3(lint_ADDR_int[5]),.T2I0(lint_ADDR_int[11]),.T2I1(lint_ADDR_int[4]),.T2I2(lint_ADDR_int[3]),.T2I3(GND),.TB2S(GND),.B2Z(NET_103),.C2Z(NET_88),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_H15_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(fpgaio_out_dup_0[25]),.T3I1(NET_37),.T3I2(NET_60),.T3I3(cnt4[0]),.TB3S(GND),.C3Z(NET_509),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_H16_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000001),.B0I0(GND),.B0I1(RESET_int[2]),.B0I2(GND),.B0I3(GND),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_in_int[68]),.T0I1(NET_36),.T0I2(NET_37),.T0I3(m0_m0_outsel_dup_0[4]),.TB0S(GND),.B0Z(not_RESET_2),.C0Z(NET_672),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H16_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_644),.T1I1(lint_ADDR_int[6]),.T1I2(NET_68),.T1I3(lint_ADDR_int[4]),.TB1S(GND),.C1Z(nx53524z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_H16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_26),.B2I1(NET_25),.B2I2(NET_23),.B2I3(NET_24),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.QST(GND),.B2Z(NET_27),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H16_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF),.QST(GND),.T3I0(NET_65),.T3I1(lint_ADDR_int[6]),.T3I2(lint_ADDR_int[2]),.T3I3(GND),.TB3S(GND),.C3Z(NET_602),.Q3Z(m0_oper1_wmode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_H17_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_36),.B0I1(fpgaio_in_int[74]),.B0I2(NET_37),.B0I3(m0_m0_control[10]),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(NET_13),.T0I1(fpgaio_out_dup_0[65]),.T0I2(NET_12),.T0I3(tcdm_result_p0[1]),.TB0S(GND),.B0Z(NET_180),.C0Z(NET_3),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(m0_m0_control[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m0_m0_control[9]),.B2I1(NET_36),.B2I2(fpgaio_in_int[73]),.B2I3(NET_37),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B2Z(NET_157),.Q2Z(m0_m0_control[9]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H17_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[3]),.T3I1(lint_ADDR_int[4]),.T3I2(lint_ADDR_int[5]),.T3I3(lint_ADDR_int[6]),.C3Z(NET_31),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H18_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_out_dup_0[33]),.B0I1(NET_6),.B0I2(NET_5),.B0I3(tcdm_rdata_p2_int[1]),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(NET_12),.T0I1(NET_13),.T0I2(fpgaio_out_dup_0[77]),.T0I3(tcdm_result_p0[13]),.TB0S(GND),.B0Z(NET_2),.C0Z(NET_237),.Q0Z(fpgaio_out_dup_0[74]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[69]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_3),.B2I1(NET_1),.B2I2(NET_2),.B2I3(NET_0),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B2Z(NET_4),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H18_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(NET_5),.T3I1(m0_m0_dataout_int[25]),.T3I2(fpgaio_out_dup_0[57]),.T3I3(NET_59),.TB3S(GND),.C3Z(NET_501),.Q3Z(fpgaio_out_dup_0[68]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_H19_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(m0_ram_control[19]),.T0I1(NET_94_CAND3_BLSTL_8_tpGCLKBUF),.T0I2(NET_103),.T0I3(m1_m0_dataout_int[19]),.TB0S(GND),.C0Z(NET_374),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx4939z1_CAND5_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[56]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H19_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B2I0(tcdm_rdata_p2_int[13]),.B2I1(NET_6),.B2I2(fpgaio_out_dup_0[45]),.B2I3(NET_5),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_out_dup_0[52]),.T2I1(NET_5),.T2I2(NET_59),.T2I3(m0_m0_dataout_int[20]),.TB2S(GND),.B2Z(NET_236),.C2Z(NET_391),.Q2Z(m0_ram_control[19]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_H19_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(NET_236),.T3I1(NET_234),.T3I2(NET_237),.T3I3(NET_235),.TB3S(GND),.C3Z(NET_238),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_H20_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(NET_94_CAND3_BLSTL_8_tpGCLKBUF),.T0I1(m1_m0_dataout_int[24]),.T0I2(m0_ram_control[24]),.T0I3(NET_103),.TB0S(GND),.C0Z(NET_484),.Q0Z(m0_ram_control[29]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H20_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[23]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_94_CAND3_BLSTL_8_tpGCLKBUF),.T1I1(m0_ram_control[23]),.T1I2(NET_103),.T1I3(m1_m0_dataout_int[23]),.TB1S(GND),.C1Z(NET_445),.Q1Z(m0_ram_control[23]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_H20_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_m0_dataout_int[22]),.B2I1(NET_94_CAND3_BLSTL_8_tpGCLKBUF),.B2I2(m0_ram_control[22]),.B2I3(NET_103),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T2I0(NET_94_CAND3_BLSTL_8_tpGCLKBUF),.T2I1(m1_m0_dataout_int[29]),.T2I2(NET_103),.T2I3(m0_ram_control[29]),.TB2S(GND),.B2Z(NET_427),.C2Z(NET_573),.Q2Z(m0_ram_control[22]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_H20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[24]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q3Z(m0_ram_control[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_28),.B0I1(fpgaio_oe_dup_0[41]),.B0I2(m1_m1_control[9]),.B0I3(NET_29_CAND4_BLSTL_8_tpGCLKBUF),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0Z(NET_159),.Q0Z(m0_ram_control[18]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[9]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_control[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H21_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T2I0(m1_m0_dataout_int[18]),.T2I1(NET_103),.T2I2(NET_94_CAND3_BLSTL_8_tpGCLKBUF),.T2I3(m0_ram_control[18]),.TB2S(GND),.C2Z(NET_355),.Q2Z(m0_ram_control[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_H21_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx4939z1_CAND5_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(m0_ram_control[17]),.T3I1(NET_103),.T3I2(m1_m0_dataout_int[17]),.T3I3(NET_94_CAND3_BLSTL_8_tpGCLKBUF),.TB3S(GND),.C3Z(NET_337),.Q3Z(fpgaio_out_dup_0[53]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_H22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx4939z1_CAND5_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[48]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H22_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_oe_dup_0[35]),.T3I1(NET_29_CAND4_BLSTL_8_tpGCLKBUF),.T3I2(m1_m1_control[3]),.T3I3(NET_28),.TB3S(GND),.C3Z(NET_693),.Q3Z(m1_m1_control[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_H23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx4939z1_CAND5_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[33]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H23_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_oe_dup_0[33]),.T3I1(NET_28),.T3I2(m1_m1_control[1]),.T3I3(NET_29_CAND4_BLSTL_8_tpGCLKBUF),.C3Z(NET_25),.Q3Z(m1_m1_control[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx4939z1_CAND5_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[36]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx4939z1_CAND5_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[42]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_tc_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_outsel_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I2_0 (.tFragBitInfo(16'b1111111100001111),.bFragBitInfo(16'b1110111000001111),.B0I0(lint_ADDR_int[14]),.B0I1(lint_ADDR_int[13]),.B0I2(lint_ADDR_int[11]),.B0I3(apb_fsm[0]),.T0I0(lint_ADDR_int[14]),.T0I1(lint_ADDR_int[13]),.T0I2(lint_ADDR_int[11]),.T0I3(apb_fsm[0]),.TB0S(m0_oper0_rdata_int[4]),.C0Z(NET_680),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_I2_1 (.tFragBitInfo(16'b1111111100001111),.bFragBitInfo(16'b1101110111010001),.B1I0(lint_ADDR_int[11]),.B1I1(apb_fsm[0]),.B1I2(lint_ADDR_int[14]),.B1I3(lint_ADDR_int[13]),.T1I0(lint_ADDR_int[14]),.T1I1(lint_ADDR_int[13]),.T1I2(lint_ADDR_int[11]),.T1I3(apb_fsm[0]),.TB1S(m0_oper0_rdata_int[5]),.C1Z(NET_660),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_I2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m0_oper1_rdata_int[3]),.B2I1(NET_45_CAND5_TLSTR_9_tpGCLKBUF),.B2I2(NET_46_CAND3_TLSTR_9_tpGCLKBUF),.B2I3(m1_oper0_rdata_int[3]),.T2I0(m0_oper1_rdata_int[3]),.T2I1(NET_45_CAND5_TLSTR_9_tpGCLKBUF),.T2I2(NET_46_CAND3_TLSTR_9_tpGCLKBUF),.T2I3(m1_oper0_rdata_int[3]),.TB2S(NET_699),.C2Z(NET_697),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_I2_3 (.tFragBitInfo(16'b1111111100001111),.bFragBitInfo(16'b1101110111010001),.B3I0(lint_ADDR_int[11]),.B3I1(apb_fsm[0]),.B3I2(lint_ADDR_int[14]),.B3I3(lint_ADDR_int[13]),.T3I0(lint_ADDR_int[14]),.T3I1(lint_ADDR_int[13]),.T3I2(lint_ADDR_int[11]),.T3I3(apb_fsm[0]),.TB3S(m0_oper0_rdata_int[3]),.C3Z(NET_699),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_I3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(m1_oper0_rdata_int[14]),.B0I1(NET_46_CAND3_TLSTR_9_tpGCLKBUF),.B0I2(m0_oper1_rdata_int[14]),.B0I3(NET_45_CAND5_TLSTR_9_tpGCLKBUF),.T0I0(m1_oper0_rdata_int[14]),.T0I1(NET_46_CAND3_TLSTR_9_tpGCLKBUF),.T0I2(m0_oper1_rdata_int[14]),.T0I3(NET_45_CAND5_TLSTR_9_tpGCLKBUF),.TB0S(NET_267),.C0Z(NET_265),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_I3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(NET_46_CAND3_TLSTR_9_tpGCLKBUF),.B1I1(m0_oper1_rdata_int[11]),.B1I2(m1_oper0_rdata_int[11]),.B1I3(NET_45_CAND5_TLSTR_9_tpGCLKBUF),.T1I0(m1_oper0_rdata_int[11]),.T1I1(NET_45_CAND5_TLSTR_9_tpGCLKBUF),.T1I2(NET_46_CAND3_TLSTR_9_tpGCLKBUF),.T1I3(m0_oper1_rdata_int[11]),.TB1S(NET_207),.C1Z(NET_205),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_I3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(m1_oper0_rdata_int[13]),.B2I1(NET_46_CAND3_TLSTR_9_tpGCLKBUF),.B2I2(m0_oper1_rdata_int[13]),.B2I3(NET_45_CAND5_TLSTR_9_tpGCLKBUF),.T2I0(m1_oper0_rdata_int[13]),.T2I1(NET_46_CAND3_TLSTR_9_tpGCLKBUF),.T2I2(m0_oper1_rdata_int[13]),.T2I3(NET_45_CAND5_TLSTR_9_tpGCLKBUF),.TB2S(NET_247),.C2Z(NET_245),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_I3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(NET_46_CAND3_TLSTR_9_tpGCLKBUF),.B3I1(NET_45_CAND5_TLSTR_9_tpGCLKBUF),.B3I2(m0_oper1_rdata_int[10]),.B3I3(m1_oper0_rdata_int[10]),.T3I0(m0_oper1_rdata_int[10]),.T3I1(m1_oper0_rdata_int[10]),.T3I2(NET_46_CAND3_TLSTR_9_tpGCLKBUF),.T3I3(NET_45_CAND5_TLSTR_9_tpGCLKBUF),.TB3S(NET_188),.C3Z(NET_186),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_I4_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B0I0(m0_m0_dataout_int[3]),.B0I1(NET_58),.B0I2(fpgaio_oe_dup_0[3]),.B0I3(NET_59),.T0I0(m0_m0_dataout_int[13]),.T0I1(NET_58),.T0I2(fpgaio_oe_dup_0[13]),.T0I3(NET_59),.TB0S(GND),.B0Z(NET_702),.C0Z(NET_250),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_I4_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(fpgaio_oe_dup_0[4]),.T1I1(NET_58),.T1I2(m0_m0_dataout_int[4]),.T1I3(NET_59),.C1Z(NET_683),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_I4_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000010),.B2I0(apb_fsm[0]),.B2I1(lint_ADDR_int[12]),.B2I2(GND),.B2I3(lint_ADDR_int[14]),.T2I0(m0_m0_dataout_int[14]),.T2I1(NET_58),.T2I2(fpgaio_oe_dup_0[14]),.T2I3(NET_59),.TB2S(GND),.B2Z(NET_46),.C2Z(NET_270),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_I4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I7_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m0_coef_wdsel_dup_0),.B0I1(NET_61),.B0I2(NET_60),.B0I3(fpgaio_out_dup_0[14]),.T0I0(NET_681),.T0I1(NET_684),.T0I2(NET_683),.T0I3(NET_682),.TB0S(GND),.B0Z(NET_271),.C0Z(NET_685),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_I7_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_270),.T1I1(NET_268),.T1I2(NET_269),.T1I3(NET_271),.C1Z(NET_272),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_I7_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.T2I0(m0_oper1_rmode_dup_0[0]),.T2I1(NET_61),.T2I2(NET_60),.T2I3(fpgaio_out_dup_0[4]),.TB2S(GND),.C2Z(NET_684),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_I7_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_703),.T3I1(NET_700),.T3I2(NET_701),.T3I3(NET_702),.TB3S(GND),.C3Z(NET_704),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_I9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_112),.B0I1(m0_m1_outsel_dup_0[2]),.B0I2(fpgaio_in_int[2]),.B0I3(NET_111),.B0Z(NET_717),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I9_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_112),.T1I1(m0_m1_tc_dup_0),.T1I2(NET_111),.T1I3(fpgaio_in_int[6]),.TB1S(GND),.C1Z(NET_635),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_I9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_112),.B2I1(m0_m1_outsel_dup_0[0]),.B2I2(fpgaio_in_int[0]),.B2I3(NET_111),.B2Z(NET_107),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I10_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(fpgaio_in_int[12]),.T1I1(NET_111),.T1I2(m0_m1_mode_dup_0[0]),.T1I3(NET_112),.C1Z(NET_225),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_I10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_467),.B2I1(NET_466),.B2I2(NET_468),.B2I3(NET_469),.B2Z(NET_458),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I10_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(fpgaio_in_int[7]),.T3I1(NET_111),.T3I2(m0_m1_control[7]),.T3I3(NET_112),.TB3S(GND),.C3Z(NET_469),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_I11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_224),.B0I1(NET_223),.B0I2(NET_222),.B0I3(NET_225),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.B0Z(NET_214),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I11_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[21]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_633),.T1I1(NET_634),.T1I2(NET_632),.T1I3(NET_635),.TB1S(GND),.C1Z(NET_624),.Q1Z(m0_m0_control[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_I11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_107),.B2I1(NET_104),.B2I2(NET_105),.B2I3(NET_106),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.B2Z(NET_79),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_control[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I12_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_679),.B0I1(NET_676),.B0I2(NET_671),.B0I3(NET_759),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.T0I0(NET_679),.T0I1(NET_676),.T0I2(NET_671),.T0I3(NET_759),.TB0S(NET_685),.Q0Z(lint_RDATA_dup_0[4]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I12_1 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.T1I0(NET_333),.T1I1(NET_332),.T1I2(NET_331),.T1I3(NET_330),.TB1S(GND),.Q1Z(lint_RDATA_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_I12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000010000000),.B2I0(NET_338),.B2I1(NET_337),.B2I2(NET_336),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.B2Z(NET_333),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I12_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.T3I0(NET_350),.T3I1(NET_352),.T3I2(NET_351),.T3I3(NET_349),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_I13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100000000000),.B0I0(NET_354),.B0I1(NET_356),.B0I2(GND),.B0I3(NET_355),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.B0Z(NET_352),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I13_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B1I0(NET_741),.B1I1(NET_304),.B1I2(NET_296),.B1I3(NET_301),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.T1I0(NET_296),.T1I1(NET_301),.T1I2(NET_741),.T1I3(NET_304),.TB1S(NET_310),.Q1Z(lint_RDATA_dup_0[15]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_I13_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_263),.B2I1(NET_258),.B2I2(NET_737),.B2I3(NET_266),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.T2I0(NET_263),.T2I1(NET_258),.T2I2(NET_737),.T2I3(NET_266),.TB2S(NET_272),.Q2Z(lint_RDATA_dup_0[14]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_I13_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.T3I0(NET_717),.T3I1(NET_716),.T3I2(NET_714),.T3I3(NET_715),.TB3S(GND),.C3Z(NET_706),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_I14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_118),.B0I1(NET_108),.B0I2(m0_m0_control[21]),.B0I3(cnt2[2]),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T0I0(NET_118),.T0I1(NET_108),.T0I2(m0_m0_control[21]),.T0I3(cnt2[2]),.TB0S(NET_417),.C0Z(NET_413),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(cnt5[0]),.B1I1(NET_118),.B1I2(NET_108),.B1I3(m0_m0_control[28]),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_108),.T1I1(m0_m0_control[28]),.T1I2(cnt5[0]),.T1I3(NET_118),.TB1S(NET_563),.C1Z(NET_559),.Q1Z(m0_m0_csel_dup_0),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_I14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_108),.B2I1(cnt5[1]),.B2I2(m0_m0_control[29]),.B2I3(NET_118),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(NET_108),.T2I1(cnt5[1]),.T2I2(m0_m0_control[29]),.T2I3(NET_118),.TB2S(NET_581),.C2Z(NET_577),.Q2Z(m0_m0_control[29]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_I14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B3I0(m0_m0_control[19]),.B3I1(NET_118),.B3I2(cnt2[0]),.B3I3(NET_108),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(cnt2[0]),.T3I1(NET_108),.T3I2(m0_m0_control[19]),.T3I3(NET_118),.TB3S(NET_382),.C3Z(NET_378),.Q3Z(m0_m0_control[19]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_I15_0 (.tFragBitInfo(16'b0001010001000100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_5__CAND5_TLSBR_9_padClk),.QRT(not_RESET_2),.QST(GND),.T0I0(GND),.T0I1(cnt5[2]),.T0I2(cnt5[0]),.T0I3(cnt5[1]),.TB0S(GND),.Q0Z(cnt5[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I15_1 (.tFragBitInfo(16'b0000000100010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_5__CAND5_TLSBR_9_padClk),.QRT(not_RESET_2),.QST(GND),.T1I0(GND),.T1I1(GND),.T1I2(cnt5[0]),.T1I3(cnt5[1]),.TB1S(GND),.Q1Z(cnt5[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_I15_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000011101110111),.B2I0(cnt5[2]),.B2I1(NET_37),.B2I2(NET_60),.B2I3(fpgaio_out_dup_0[30]),.QCK(CLK_int_5__CAND5_TLSBR_9_padClk),.QRT(not_RESET_2),.QST(GND),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(RESET_int[1]),.TB2S(GND),.B2Z(NET_598),.C2Z(not_RESET_1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I15_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_5__CAND5_TLSBR_9_padClk),.QRT(not_RESET_2),.QST(GND),.T3I0(GND),.T3I1(GND),.T3I2(cnt5[0]),.T3I3(GND),.TB3S(GND),.Q3Z(cnt5[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_I16_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_675),.B0I1(NET_673),.B0I2(NET_672),.B0I3(NET_674),.QCK(CLK_int_2__CAND2_TLSBR_9_padClk),.QRT(not_RESET_2),.QST(GND),.T0I0(m0_m0_outsel_dup_0[5]),.T0I1(fpgaio_in_int[69]),.T0I2(NET_36),.T0I3(NET_37),.TB0S(GND),.B0Z(NET_676),.C0Z(NET_652),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I16_1 (.tFragBitInfo(16'b0001001100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_2__CAND2_TLSBR_9_padClk),.QRT(not_RESET_2),.QST(GND),.T1I0(cnt2[1]),.T1I1(GND),.T1I2(cnt2[0]),.T1I3(cnt2[2]),.TB1S(GND),.Q1Z(cnt2[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_I16_2 (.tFragBitInfo(16'b0000000000010010),.bFragBitInfo(16'b0000011101110111),.B2I0(fpgaio_out_dup_0[20]),.B2I1(NET_60),.B2I2(cnt2[1]),.B2I3(NET_37),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_2__CAND2_TLSBR_9_padClk),.QRT(not_RESET_2),.QST(GND),.T2I0(cnt2[1]),.T2I1(GND),.T2I2(cnt2[0]),.T2I3(GND),.TB2S(GND),.B2Z(NET_399),.Q2Z(cnt2[1]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_I16_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_2__CAND2_TLSBR_9_padClk),.QRT(not_RESET_2),.QST(GND),.T3I0(GND),.T3I1(GND),.T3I2(cnt2[0]),.T3I3(GND),.TB3S(GND),.Q3Z(cnt2[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_I17_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_259),.B0I1(NET_262),.B0I2(NET_260),.B0I3(NET_261),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T0I0(NET_297),.T0I1(NET_298),.T0I2(NET_300),.T0I3(NET_299),.TB0S(GND),.B0Z(NET_263),.C0Z(NET_301),.Q0Z(m0_m0_control[8]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I17_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_in_int[72]),.T1I1(NET_36),.T1I2(NET_37),.T1I3(m0_m0_control[8]),.C1Z(NET_278),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_I17_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B2I0(fpgaio_in_int[79]),.B2I1(NET_36),.B2I2(m0_m0_csel_dup_0),.B2I3(NET_37),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T2I0(m0_m0_mode_dup_0[1]),.T2I1(NET_36),.T2I2(NET_37),.T2I3(fpgaio_in_int[77]),.TB2S(GND),.B2Z(NET_297),.C2Z(NET_239),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I18_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_667),.B0I1(NET_668),.B0I2(NET_670),.B0I3(NET_669),.T0I0(NET_6),.T0I1(fpgaio_out_dup_0[36]),.T0I2(NET_5),.T0I3(tcdm_rdata_p2_int[4]),.TB0S(GND),.B0Z(NET_671),.C0Z(NET_669),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_I18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I18_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_13),.B2I1(fpgaio_out_dup_0[79]),.B2I2(tcdm_result_p0[15]),.B2I3(NET_12),.T2I0(fpgaio_out_dup_0[78]),.T2I1(tcdm_result_p0[14]),.T2I2(NET_12),.T2I3(NET_13),.TB2S(GND),.B2Z(NET_295),.C2Z(NET_257),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_I18_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_13),.T3I1(tcdm_result_p0[4]),.T3I2(NET_12),.T3I3(fpgaio_out_dup_0[68]),.TB3S(GND),.C3Z(NET_670),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_I19_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_out_dup_0[46]),.B0I1(tcdm_rdata_p2_int[14]),.B0I2(NET_5),.B0I3(NET_6),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_out_dup_0[47]),.T0I1(NET_5),.T0I2(tcdm_rdata_p2_int[15]),.T0I3(NET_6),.TB0S(GND),.B0Z(NET_256),.C0Z(NET_294),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I19_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[48]),.T1I1(NET_59),.T1I2(NET_5),.T1I3(m0_m0_dataout_int[16]),.TB1S(GND),.C1Z(NET_317),.Q1Z(m0_coef_wdsel_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_I19_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_294),.B2I1(NET_292),.B2I2(NET_295),.B2I3(NET_293),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T2I0(NET_255),.T2I1(NET_254),.T2I2(NET_257),.T2I3(NET_256),.TB2S(GND),.B2Z(NET_296),.C2Z(NET_258),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q0Z(m0_ram_control[25]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_control[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_m0_dataout_int[25]),.B2I1(m0_ram_control[25]),.B2I2(NET_18_CAND4_BLSTR_9_tpGCLKBUF),.B2I3(NET_61),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2Z(NET_510),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I20_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_oe_dup_0[42]),.T3I1(NET_29),.T3I2(m1_m1_control[10]),.T3I3(NET_28_CAND5_BLSTR_9_tpGCLKBUF),.TB3S(GND),.C3Z(NET_182),.Q3Z(fpgaio_out_dup_0[58]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_I21_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx49871z1_CAND3_BLSTR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T0I0(NET_17_CAND2_BLSTR_9_tpGCLKBUF),.T0I1(m1_m0_dataout_int[15]),.T0I2(NET_18_CAND4_BLSTR_9_tpGCLKBUF),.T0I3(m1_ram_control[15]),.TB0S(GND),.C0Z(NET_293),.Q0Z(m1_ram_control[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I21_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx49871z1_CAND3_BLSTR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(m1_ram_control[13]),.T1I1(NET_17_CAND2_BLSTR_9_tpGCLKBUF),.T1I2(NET_18_CAND4_BLSTR_9_tpGCLKBUF),.T1I3(m1_m0_dataout_int[13]),.C1Z(NET_235),.Q1Z(m1_ram_control[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_I21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_17_CAND2_BLSTR_9_tpGCLKBUF),.B2I1(m1_m0_dataout_int[14]),.B2I2(NET_18_CAND4_BLSTR_9_tpGCLKBUF),.B2I3(m1_ram_control[14]),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx49871z1_CAND3_BLSTR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2Z(NET_255),.Q2Z(m1_ram_control[13]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I21_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx49871z1_CAND3_BLSTR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_17_CAND2_BLSTR_9_tpGCLKBUF),.T3I1(m1_ram_control[4]),.T3I2(NET_18_CAND4_BLSTR_9_tpGCLKBUF),.T3I3(m1_m0_dataout_int[4]),.C3Z(NET_668),.Q3Z(m1_ram_control[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_I23_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_28_CAND5_BLSTR_9_tpGCLKBUF),.B0I1(fpgaio_oe_dup_0[47]),.B0I2(m1_m1_csel_dup_0),.B0I3(NET_29),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T0I0(NET_29),.T0I1(NET_28_CAND5_BLSTR_9_tpGCLKBUF),.T0I2(m1_m1_mode_dup_0[1]),.T0I3(fpgaio_oe_dup_0[45]),.TB0S(GND),.B0Z(NET_299),.C0Z(NET_241),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I23_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_osel_dup_0),.T1I1(NET_28_CAND5_BLSTR_9_tpGCLKBUF),.T1I2(fpgaio_oe_dup_0[46]),.T1I3(NET_29),.TB1S(GND),.C1Z(NET_261),.Q1Z(m1_m1_csel_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_I23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_mode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[46]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[55]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_outsel_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_outsel_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.Q3Z(m1_m0_outsel_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I31_2 (.tFragBitInfo(16'b1010101011111111),.bFragBitInfo(16'b1010100011111101),.B2I0(apb_fsm[0]),.B2I1(lint_ADDR_int[12]),.B2I2(lint_ADDR_int[13]),.B2I3(lint_ADDR_int[11]),.T2I0(apb_fsm[0]),.T2I1(lint_ADDR_int[12]),.T2I2(lint_ADDR_int[13]),.T2I3(lint_ADDR_int[11]),.TB2S(m1_oper0_rdata_int[31]),.C2Z(NET_752),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_I31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I32_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m1_oper0_rdata_int[22]),.T1I1(m1_coef_rdata_int[22]),.T1I2(NET_45_CAND5_BLSBR_9_tpGCLKBUF),.T1I3(NET_43_CAND3_BLSBR_9_tpGCLKBUF),.C1Z(NET_436),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_I32_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_45_CAND5_BLSBR_9_tpGCLKBUF),.B2I1(NET_43_CAND3_BLSBR_9_tpGCLKBUF),.B2I2(m1_oper0_rdata_int[28]),.B2I3(m1_coef_rdata_int[28]),.T2I0(m1_coef_rdata_int[21]),.T2I1(m1_oper0_rdata_int[21]),.T2I2(NET_43_CAND3_BLSBR_9_tpGCLKBUF),.T2I3(NET_45_CAND5_BLSBR_9_tpGCLKBUF),.TB2S(GND),.B2Z(NET_564),.C2Z(NET_418),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_I32_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m1_oper0_rdata_int[29]),.T3I1(NET_45_CAND5_BLSBR_9_tpGCLKBUF),.T3I2(NET_43_CAND3_BLSBR_9_tpGCLKBUF),.T3I3(m1_coef_rdata_int[29]),.C3Z(NET_582),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J1_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.T0I0(NET_117),.T0I1(NET_46_CAND3_TLSTR_10_tpGCLKBUF),.T0I2(m0_oper1_rdata_int[12]),.T0I3(m0_oper0_rdata_int[12]),.TB0S(GND),.C0Z(NET_227),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J1_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_41_CAND4_TLSTR_10_tpGCLKBUF),.T2I1(m0_coef_rdata_int[29]),.T2I2(NET_46_CAND3_TLSTR_10_tpGCLKBUF),.T2I3(m0_oper1_rdata_int[29]),.TB2S(GND),.C2Z(NET_584),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J1_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m0_oper1_rdata_int[7]),.T3I1(m0_oper0_rdata_int[7]),.T3I2(NET_46_CAND3_TLSTR_10_tpGCLKBUF),.T3I3(NET_117),.TB3S(GND),.C3Z(NET_471),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J2_0 (.tFragBitInfo(16'b0010101000000000),.bFragBitInfo(16'b0000100010001000),.B0I0(NET_658),.B0I1(NET_657),.B0I2(NET_41_CAND4_TLSTR_10_tpGCLKBUF),.B0I3(m0_coef_rdata_int[5]),.T0I0(NET_696),.T0I1(m0_coef_rdata_int[3]),.T0I2(NET_41_CAND4_TLSTR_10_tpGCLKBUF),.T0I3(NET_697),.TB0S(GND),.B0Z(NET_659),.C0Z(NET_698),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(NET_46_CAND3_TLSTR_10_tpGCLKBUF),.B1I1(m0_oper1_rdata_int[15]),.B1I2(m1_oper0_rdata_int[15]),.B1I3(NET_45_CAND5_TLSTR_10_tpGCLKBUF),.T1I0(m1_oper0_rdata_int[15]),.T1I1(NET_45_CAND5_TLSTR_10_tpGCLKBUF),.T1I2(NET_46_CAND3_TLSTR_10_tpGCLKBUF),.T1I3(m0_oper1_rdata_int[15]),.TB1S(NET_305),.C1Z(NET_303),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_J2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_45_CAND5_TLSTR_10_tpGCLKBUF),.B2I1(m0_oper1_rdata_int[5]),.B2I2(NET_46_CAND3_TLSTR_10_tpGCLKBUF),.B2I3(m1_oper0_rdata_int[5]),.T2I0(NET_45_CAND5_TLSTR_10_tpGCLKBUF),.T2I1(m0_oper1_rdata_int[5]),.T2I2(NET_46_CAND3_TLSTR_10_tpGCLKBUF),.T2I3(m1_oper0_rdata_int[5]),.TB2S(NET_660),.C2Z(NET_658),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B3I0(m0_oper1_rdata_int[8]),.B3I1(NET_46_CAND3_TLSTR_10_tpGCLKBUF),.B3I2(m1_oper0_rdata_int[8]),.B3I3(NET_45_CAND5_TLSTR_10_tpGCLKBUF),.T3I0(m1_oper0_rdata_int[8]),.T3I1(NET_45_CAND5_TLSTR_10_tpGCLKBUF),.T3I2(m0_oper1_rdata_int[8]),.T3I3(NET_46_CAND3_TLSTR_10_tpGCLKBUF),.TB3S(NET_286),.C3Z(NET_284),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J3_0 (.tFragBitInfo(16'b0010101000000000),.bFragBitInfo(16'b0000100010001000),.B0I0(NET_264),.B0I1(NET_265),.B0I2(m0_coef_rdata_int[14]),.B0I3(NET_41_CAND4_TLSTR_10_tpGCLKBUF),.T0I0(NET_303),.T0I1(m0_coef_rdata_int[15]),.T0I2(NET_41_CAND4_TLSTR_10_tpGCLKBUF),.T0I3(NET_302),.TB0S(GND),.B0Z(NET_266),.C0Z(NET_304),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J3_1 (.tFragBitInfo(16'b0010101000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_283),.T1I1(m0_coef_rdata_int[8]),.T1I2(NET_41_CAND4_TLSTR_10_tpGCLKBUF),.T1I3(NET_284),.TB1S(GND),.C1Z(NET_285),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_J3_2 (.tFragBitInfo(16'b0100110000000000),.bFragBitInfo(16'b0010101000000000),.B2I0(NET_245),.B2I1(m0_coef_rdata_int[13]),.B2I2(NET_41_CAND4_TLSTR_10_tpGCLKBUF),.B2I3(NET_244),.T2I0(m0_coef_rdata_int[10]),.T2I1(NET_186),.T2I2(NET_41_CAND4_TLSTR_10_tpGCLKBUF),.T2I3(NET_185),.TB2S(GND),.B2Z(NET_246),.C2Z(NET_187),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J3_3 (.tFragBitInfo(16'b0000100010001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_204),.T3I1(NET_205),.T3I2(m0_coef_rdata_int[11]),.T3I3(NET_41_CAND4_TLSTR_10_tpGCLKBUF),.TB3S(GND),.C3Z(NET_206),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J4_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_58),.B0I1(m0_m0_dataout_int[9]),.B0I2(fpgaio_oe_dup_0[9]),.B0I3(NET_59),.T0I0(NET_59),.T0I1(NET_58),.T0I2(fpgaio_oe_dup_0[11]),.T0I3(m0_m0_dataout_int[11]),.TB0S(GND),.B0Z(NET_168),.C0Z(NET_210),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J4_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(fpgaio_oe_dup_0[8]),.T1I1(NET_58),.T1I2(m0_m0_dataout_int[8]),.T1I3(NET_59),.C1Z(NET_289),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J4_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_58),.T2I1(fpgaio_oe_dup_0[10]),.T2I2(NET_59),.T2I3(m0_m0_dataout_int[10]),.TB2S(GND),.C2Z(NET_191),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J4_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m0_m0_dataout_int[5]),.T3I1(NET_58),.T3I2(NET_59),.T3I3(fpgaio_oe_dup_0[5]),.C3Z(NET_663),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000100),.B2I0(lint_ADDR_int[14]),.B2I1(apb_fsm[0]),.B2I2(lint_ADDR_int[13]),.B2I3(GND),.B2Z(NET_117),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J7_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B0I0(fpgaio_out_dup_0[13]),.B0I1(NET_60),.B0I2(m0_oper1_wdsel_dup_0),.B0I3(NET_61),.T0I0(m0_oper1_rmode_dup_0[1]),.T0I1(NET_60),.T0I2(NET_61),.T0I3(fpgaio_out_dup_0[5]),.TB0S(GND),.B0Z(NET_251),.C0Z(NET_664),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J7_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_663),.T1I1(NET_664),.T1I2(NET_661),.T1I3(NET_662),.TB1S(GND),.C1Z(NET_665),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_J7_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_250),.B2I1(NET_248),.B2I2(NET_251),.B2I3(NET_249),.T2I0(fpgaio_out_dup_0[8]),.T2I1(NET_60),.T2I2(NET_61),.T2I3(m0_coef_rmode_dup_0[0]),.TB2S(GND),.B2Z(NET_252),.C2Z(NET_290),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J8_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_189),.B0I1(NET_192),.B0I2(NET_191),.B0I3(NET_190),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.T0I0(NET_167),.T0I1(NET_168),.T0I2(NET_169),.T0I3(NET_166),.TB0S(GND),.B0Z(NET_193),.C0Z(NET_170),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.Q1Z(m0_m0_rnd_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J8_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_60),.B2I1(m0_coef_wmode_dup_0[0]),.B2I2(fpgaio_out_dup_0[10]),.B2I3(NET_61),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.T2I0(NET_60),.T2I1(m0_coef_rmode_dup_0[1]),.T2I2(NET_61),.T2I3(fpgaio_out_dup_0[9]),.TB2S(GND),.B2Z(NET_192),.C2Z(NET_169),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J9_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_473),.B0I1(NET_470),.B0I2(NET_471),.B0I3(NET_472),.T0I0(NET_290),.T0I1(NET_289),.T0I2(NET_288),.T0I3(NET_287),.TB0S(GND),.B0Z(NET_467),.C0Z(NET_291),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J9_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_41),.T1I1(NET_43),.T1I2(m1_coef_rdata_int[12]),.T1I3(m0_coef_rdata_int[12]),.TB1S(GND),.C1Z(NET_228),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_J9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_227),.B2I1(NET_226),.B2I2(NET_228),.B2I3(NET_229),.B2Z(NET_223),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J9_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_41),.T3I1(NET_43),.T3I2(m0_coef_rdata_int[7]),.T3I3(m1_coef_rdata_int[7]),.TB3S(GND),.C3Z(NET_472),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_rmode_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J10_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_209),.T1I1(NET_208),.T1I2(NET_211),.T1I3(NET_210),.C1Z(NET_212),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J10_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_61),.T3I1(NET_60),.T3I2(fpgaio_out_dup_0[11]),.T3I3(m0_coef_wmode_dup_0[1]),.C3Z(NET_211),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J11_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T0I0(NET_44),.T0I1(m1_oper1_rdata_int[29]),.T0I2(m0_oper0_rdata_int[29]),.T0I3(NET_117),.TB0S(GND),.C0Z(NET_583),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J11_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_44),.T1I1(m1_oper1_rdata_int[28]),.T1I2(m0_oper0_rdata_int[28]),.T1I3(NET_117),.TB1S(GND),.C1Z(NET_565),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_J11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010101000000000),.B2I0(NET_564),.B2I1(tcdm_rdata_p0_int[28]),.B2I2(NET_124),.B2I3(NET_565),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T2I0(NET_564),.T2I1(tcdm_rdata_p0_int[28]),.T2I2(NET_124),.T2I3(NET_565),.TB2S(NET_566),.C2Z(NET_549),.Q2Z(m0_m0_mode_dup_0[1]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_J11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000011000000),.B3I0(NET_124),.B3I1(NET_582),.B3I2(NET_583),.B3I3(tcdm_rdata_p0_int[29]),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_583),.T3I1(tcdm_rdata_p0_int[29]),.T3I2(NET_124),.T3I3(NET_582),.TB3S(NET_584),.C3Z(NET_567),.Q3Z(m0_coef_rmode_dup_0[1]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_J12_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_690),.B0I1(NET_698),.B0I2(NET_761),.B0I3(NET_695),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T0I0(NET_690),.T0I1(NET_698),.T0I2(NET_761),.T0I3(NET_695),.TB0S(NET_704),.Q0Z(lint_RDATA_dup_0[3]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J12_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_659),.B2I1(NET_656),.B2I2(NET_757),.B2I3(NET_651),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T2I0(NET_659),.T2I1(NET_656),.T2I2(NET_757),.T2I3(NET_651),.TB2S(NET_665),.Q2Z(lint_RDATA_dup_0[5]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_J12_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_246),.B3I1(NET_735),.B3I2(NET_243),.B3I3(NET_238),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T3I0(NET_243),.T3I1(NET_238),.T3I2(NET_246),.T3I3(NET_735),.TB3S(NET_252),.Q3Z(lint_RDATA_dup_0[13]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_J13_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_198),.B0I1(NET_206),.B0I2(NET_203),.B0I3(NET_733),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T0I0(NET_198),.T0I1(NET_206),.T0I2(NET_203),.T0I3(NET_733),.TB0S(NET_212),.Q0Z(lint_RDATA_dup_0[11]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B1I0(fpgaio_out_dup_0[50]),.B1I1(tcdm_result_p3[18]),.B1I2(NET_96),.B1I3(NET_99),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T1I0(NET_96),.T1I1(NET_99),.T1I2(fpgaio_out_dup_0[50]),.T1I3(tcdm_result_p3[18]),.TB1S(NET_357),.C1Z(NET_354),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_J13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_96),.B2I1(fpgaio_out_dup_0[56]),.B2I2(tcdm_result_p3[24]),.B2I3(NET_99),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T2I0(NET_96),.T2I1(fpgaio_out_dup_0[56]),.T2I2(tcdm_result_p3[24]),.T2I3(NET_99),.TB2S(NET_486),.C2Z(NET_483),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J13_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_179),.B3I1(NET_184),.B3I2(NET_731),.B3I3(NET_187),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T3I0(NET_731),.T3I1(NET_187),.T3I2(NET_179),.T3I3(NET_184),.TB3S(NET_193),.Q3Z(lint_RDATA_dup_0[10]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_J14_0 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000000000100),.B0I0(GND),.B0I1(lint_ADDR_int[6]),.B0I2(lint_ADDR_int[5]),.B0I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T0I0(apb_fsm[0]),.T0I1(lint_ADDR_int[13]),.T0I2(lint_ADDR_int[14]),.T0I3(GND),.TB0S(GND),.B0Z(NET_9),.C0Z(NET_43),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(tcdm_result_p3[21]),.B1I1(NET_99),.B1I2(fpgaio_out_dup_0[53]),.B1I3(NET_96),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T1I0(fpgaio_out_dup_0[53]),.T1I1(NET_96),.T1I2(tcdm_result_p3[21]),.T1I3(NET_99),.TB1S(NET_411),.C1Z(NET_408),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_J14_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_277),.B2I1(NET_282),.B2I2(NET_285),.B2I3(NET_739),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T2I0(NET_277),.T2I1(NET_282),.T2I2(NET_285),.T2I3(NET_739),.TB2S(NET_291),.Q2Z(lint_RDATA_dup_0[8]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_J14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B3I0(tcdm_result_p3[26]),.B3I1(NET_99),.B3I2(fpgaio_out_dup_0[58]),.B3I3(NET_96),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T3I0(fpgaio_out_dup_0[58]),.T3I1(NET_96),.T3I2(tcdm_result_p3[26]),.T3I3(NET_99),.TB3S(NET_521),.C3Z(NET_518),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_J15_0 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000000000010000),.B0I0(lint_ADDR_int[15]),.B0I1(lint_ADDR_int[14]),.B0I2(NET_73),.B0I3(lint_ADDR_int[12]),.T0I0(NET_73),.T0I1(NET_71),.T0I2(GND),.T0I3(NET_72),.TB0S(GND),.B0Z(NET_149),.C0Z(NET_69),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(tcdm_result_p3[19]),.B1I1(NET_99),.B1I2(fpgaio_out_dup_0[51]),.B1I3(NET_96),.T1I0(fpgaio_out_dup_0[51]),.T1I1(NET_96),.T1I2(tcdm_result_p3[19]),.T1I3(NET_99),.TB1S(NET_376),.C1Z(NET_373),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_J15_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000001000000),.B2I0(lint_ADDR_int[15]),.B2I1(lint_ADDR_int[14]),.B2I2(NET_73),.B2I3(lint_ADDR_int[12]),.T2I0(GND),.T2I1(lint_ADDR_int[14]),.T2I2(lint_ADDR_int[13]),.T2I3(lint_ADDR_int[12]),.TB2S(GND),.B2Z(NET_171),.C2Z(NET_74),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J15_3 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int[15]),.T3I1(lint_ADDR_int[8]),.T3I2(NET_74),.T3I3(lint_ADDR_int[10]),.C3Z(NET_72),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J16_0 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_652),.B0I1(NET_653),.B0I2(NET_655),.B0I3(NET_654),.T0I0(NET_8),.T0I1(NET_11),.T0I2(NET_9),.T0I3(GND),.TB0S(GND),.B0Z(NET_656),.C0Z(NET_60),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J16_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_200),.T1I1(NET_199),.T1I2(NET_201),.T1I3(NET_202),.C1Z(NET_203),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_602),.B2I1(NET_69),.B2I2(NET_148),.B2I3(NET_70),.B2Z(nx4939z1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J16_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_693),.T3I1(NET_692),.T3I2(NET_691),.T3I3(NET_694),.C3Z(NET_695),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J17_0 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_239),.B0I1(NET_240),.B0I2(NET_241),.B0I3(NET_242),.T0I0(NET_31),.T0I1(NET_8),.T0I2(GND),.T0I3(GND),.TB0S(GND),.B0Z(NET_243),.C0Z(NET_32),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J17_2 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_182),.B2I1(NET_180),.B2I2(NET_183),.B2I3(NET_181),.T2I0(GND),.T2I1(NET_11),.T2I2(NET_10),.T2I3(NET_9),.TB2S(GND),.B2Z(NET_184),.C2Z(NET_5),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J17_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_278),.T3I1(NET_281),.T3I2(NET_280),.T3I3(NET_279),.TB3S(GND),.C3Z(NET_282),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J18_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_13),.B0I1(tcdm_result_p0[8]),.B0I2(fpgaio_out_dup_0[72]),.B0I3(NET_12),.T0I0(NET_13),.T0I1(tcdm_result_p0[10]),.T0I2(fpgaio_out_dup_0[74]),.T0I3(NET_12),.TB0S(GND),.B0Z(NET_276),.C0Z(NET_178),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J18_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_274),.T1I1(NET_276),.T1I2(NET_273),.T1I3(NET_275),.C1Z(NET_277),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J18_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_5),.B2I1(fpgaio_out_dup_0[42]),.B2I2(tcdm_rdata_p2_int[10]),.B2I3(NET_6),.T2I0(NET_175),.T2I1(NET_176),.T2I2(NET_177),.T2I3(NET_178),.TB2S(GND),.B2Z(NET_177),.C2Z(NET_179),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J18_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_13),.T3I1(tcdm_result_p0[11]),.T3I2(NET_12),.T3I3(fpgaio_out_dup_0[75]),.TB3S(GND),.C3Z(NET_197),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_317),.B0I1(NET_319),.B0I2(NET_318),.B0I3(NET_320),.B0Z(NET_314),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J19_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_647),.T1I1(NET_650),.T1I2(NET_649),.T1I3(NET_648),.TB1S(GND),.C1Z(NET_651),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_J19_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_194),.B2I1(NET_197),.B2I2(NET_195),.B2I3(NET_196),.T2I0(NET_5),.T2I1(fpgaio_out_dup_0[37]),.T2I2(NET_6),.T2I3(tcdm_rdata_p2_int[5]),.TB2S(GND),.B2Z(NET_198),.C2Z(NET_649),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J19_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_5),.T3I1(fpgaio_out_dup_0[43]),.T3I2(tcdm_rdata_p2_int[11]),.T3I3(NET_6),.C3Z(NET_196),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J20_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx49871z1_CAND3_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T0I0(m1_m0_dataout_int[16]),.T0I1(m0_ram_control[16]),.T0I2(NET_18_CAND4_BLSTR_10_tpGCLKBUF),.T0I3(NET_61),.TB0S(GND),.C0Z(NET_327),.Q0Z(m1_ram_control[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J20_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T2I0(NET_18_CAND4_BLSTR_10_tpGCLKBUF),.T2I1(m1_m0_dataout_int[5]),.T2I2(NET_17_CAND2_BLSTR_10_tpGCLKBUF),.T2I3(m1_ram_control[5]),.TB2S(GND),.C2Z(NET_648),.Q2Z(m0_ram_control[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_J20_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx49871z1_CAND3_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_dataout_int[10]),.T3I1(NET_17_CAND2_BLSTR_10_tpGCLKBUF),.T3I2(m1_ram_control[10]),.T3I3(NET_18_CAND4_BLSTR_10_tpGCLKBUF),.C3Z(NET_176),.Q3Z(m1_ram_control[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_18_CAND4_BLSTR_10_tpGCLKBUF),.B0I1(NET_17_CAND2_BLSTR_10_tpGCLKBUF),.B0I2(m1_m0_dataout_int[11]),.B0I3(m1_ram_control[11]),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B0Z(NET_195),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[8]),.Q1EN(nx49871z1_CAND3_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q1Z(m1_ram_control[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wmode_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J21_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx49871z1_CAND3_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_18_CAND4_BLSTR_10_tpGCLKBUF),.T3I1(NET_17_CAND2_BLSTR_10_tpGCLKBUF),.T3I2(m1_ram_control[8]),.T3I3(m1_m0_dataout_int[8]),.TB3S(GND),.C3Z(NET_274),.Q3Z(m1_ram_control[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_J24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[61]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_32),.B0I1(NET_33),.B0I2(m1_m1_dataout_int[8]),.B0I3(m1_m0_control[8]),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B0Z(NET_281),.Q0Z(m1_m0_control[8]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_mode_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_32),.B0I1(m1_m1_dataout_int[16]),.B0I2(m1_m0_rnd_dup_0),.B0I3(NET_33),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B0Z(NET_318),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_rnd_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J30_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(m1_m1_dataout_int[5]),.B0I1(m1_m0_outsel_dup_0[5]),.B0I2(NET_33),.B0I3(NET_32),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T0I0(NET_32),.T0I1(m1_m1_dataout_int[3]),.T0I2(NET_33),.T0I3(m1_m0_outsel_dup_0[3]),.TB0S(GND),.B0Z(NET_655),.C0Z(NET_694),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J30_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(m1_m0_osel_dup_0),.T1I1(m1_m1_dataout_int[14]),.T1I2(NET_33),.T1I3(NET_32),.TB1S(GND),.C1Z(NET_262),.Q1Z(m1_m0_csel_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_J30_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_32),.B2I1(m1_m1_dataout_int[1]),.B2I2(NET_33),.B2I3(m1_m0_outsel_dup_0[1]),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T2I0(NET_32),.T2I1(m1_m1_dataout_int[15]),.T2I2(m1_m0_csel_dup_0),.T2I3(NET_33),.TB2S(GND),.B2Z(NET_26),.C2Z(NET_300),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J30_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_32),.T3I1(m1_m1_dataout_int[4]),.T3I2(NET_33),.T3I3(m1_m0_outsel_dup_0[4]),.TB3S(GND),.C3Z(NET_675),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_J31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_44_CAND4_BLSBR_10_tpGCLKBUF),.B0I1(m1_coef_rdata_int[3]),.B0I2(NET_43_CAND3_BLSBR_10_tpGCLKBUF),.B0I3(m1_oper1_rdata_int[3]),.B0Z(NET_696),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J31_3 (.tFragBitInfo(16'b1111111100110011),.bFragBitInfo(16'b1100100011111011),.B3I0(lint_ADDR_int[12]),.B3I1(apb_fsm[0]),.B3I2(lint_ADDR_int[13]),.B3I3(lint_ADDR_int[11]),.T3I0(lint_ADDR_int[13]),.T3I1(lint_ADDR_int[11]),.T3I2(lint_ADDR_int[12]),.T3I3(apb_fsm[0]),.TB3S(m1_oper0_rdata_int[25]),.C3Z(NET_746),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J32_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B0I0(m1_coef_rdata_int[19]),.B0I1(NET_45_CAND5_BLSBR_10_tpGCLKBUF),.B0I2(NET_43_CAND3_BLSBR_10_tpGCLKBUF),.B0I3(m1_oper0_rdata_int[19]),.T0I0(m1_coef_rdata_int[18]),.T0I1(NET_45_CAND5_BLSBR_10_tpGCLKBUF),.T0I2(NET_43_CAND3_BLSBR_10_tpGCLKBUF),.T0I3(m1_oper0_rdata_int[18]),.TB0S(GND),.B0Z(NET_383),.C0Z(NET_364),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J32_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m1_oper1_rdata_int[15]),.T1I1(m1_coef_rdata_int[15]),.T1I2(NET_43_CAND3_BLSBR_10_tpGCLKBUF),.T1I3(NET_44_CAND4_BLSBR_10_tpGCLKBUF),.C1Z(NET_302),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J32_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_44_CAND4_BLSBR_10_tpGCLKBUF),.B2I1(m1_oper0_rdata_int[12]),.B2I2(NET_45_CAND5_BLSBR_10_tpGCLKBUF),.B2I3(m1_oper1_rdata_int[12]),.T2I0(m1_coef_rdata_int[24]),.T2I1(m1_oper0_rdata_int[24]),.T2I2(NET_43_CAND3_BLSBR_10_tpGCLKBUF),.T2I3(NET_45_CAND5_BLSBR_10_tpGCLKBUF),.TB2S(GND),.B2Z(NET_229),.C2Z(NET_493),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J32_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m1_oper1_rdata_int[7]),.T3I1(m1_oper0_rdata_int[7]),.T3I2(NET_44_CAND4_BLSBR_10_tpGCLKBUF),.T3I3(NET_45_CAND5_BLSBR_10_tpGCLKBUF),.C3Z(NET_473),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_K1_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T0I0(NET_117),.T0I1(NET_46_CAND3_TLSTR_11_tpGCLKBUF),.T0I2(m0_oper1_rdata_int[2]),.T0I3(m0_oper0_rdata_int[2]),.TB0S(GND),.C0Z(NET_719),.Q0Z(m0_coef_wdata_dup_0[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K1_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_117),.T1I1(m0_oper1_rdata_int[6]),.T1I2(m0_oper0_rdata_int[6]),.T1I3(NET_46_CAND3_TLSTR_11_tpGCLKBUF),.C1Z(NET_637),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[27]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K1_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(NET_117),.T3I1(m0_oper1_rdata_int[0]),.T3I2(NET_46_CAND3_TLSTR_11_tpGCLKBUF),.T3I3(m0_oper0_rdata_int[0]),.TB3S(GND),.C3Z(NET_114),.Q3Z(m0_coef_wdata_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[29]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B1I0(NET_46_CAND3_TLSTR_11_tpGCLKBUF),.B1I1(NET_45_CAND5_TLSTR_11_tpGCLKBUF),.B1I2(m1_oper0_rdata_int[9]),.B1I3(m0_oper1_rdata_int[9]),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T1I0(m1_oper0_rdata_int[9]),.T1I1(m0_oper1_rdata_int[9]),.T1I2(NET_46_CAND3_TLSTR_11_tpGCLKBUF),.T1I3(NET_45_CAND5_TLSTR_11_tpGCLKBUF),.TB1S(NET_165),.C1Z(NET_163),.Q1Z(m0_coef_wdata_dup_0[30]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_K2_2 (.tFragBitInfo(16'b0100110000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T2I0(m0_coef_rdata_int[4]),.T2I1(NET_677),.T2I2(NET_41_CAND4_TLSTR_11_tpGCLKBUF),.T2I3(NET_678),.TB2S(GND),.C2Z(NET_679),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B3I0(m1_oper0_rdata_int[4]),.B3I1(NET_45_CAND5_TLSTR_11_tpGCLKBUF),.B3I2(m0_oper1_rdata_int[4]),.B3I3(NET_46_CAND3_TLSTR_11_tpGCLKBUF),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(m0_oper1_rdata_int[4]),.T3I1(NET_46_CAND3_TLSTR_11_tpGCLKBUF),.T3I2(m1_oper0_rdata_int[4]),.T3I3(NET_45_CAND5_TLSTR_11_tpGCLKBUF),.TB3S(NET_680),.C3Z(NET_678),.Q3Z(m0_coef_wdata_dup_0[28]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K3_0 (.tFragBitInfo(16'b0100110000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T0I0(m0_coef_rdata_int[9]),.T0I1(NET_163),.T0I2(NET_41_CAND4_TLSTR_11_tpGCLKBUF),.T0I3(NET_162),.TB0S(GND),.C0Z(NET_164),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K4_0 (.tFragBitInfo(16'b0100110000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(lint_ADDR_int[12]),.B0I1(NET_65),.B0I2(lint_ADDR_int[13]),.B0I3(NET_144),.T0I0(m0_coef_rdata_int[1]),.T0I1(NET_39),.T0I2(NET_41_CAND4_TLSTR_11_tpGCLKBUF),.T0I3(NET_40),.TB0S(GND),.B0Z(nx15998z1),.C0Z(NET_42),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B1I0(m0_oper1_rdata_int[1]),.B1I1(m1_oper0_rdata_int[1]),.B1I2(NET_45_CAND5_TLSTR_11_tpGCLKBUF),.B1I3(NET_46_CAND3_TLSTR_11_tpGCLKBUF),.T1I0(NET_45_CAND5_TLSTR_11_tpGCLKBUF),.T1I1(NET_46_CAND3_TLSTR_11_tpGCLKBUF),.T1I2(m0_oper1_rdata_int[1]),.T1I3(m1_oper0_rdata_int[1]),.TB1S(NET_47),.C1Z(NET_40),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_K4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K6_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_WEN_int),.T1I1(lint_ADDR_int[14]),.T1I2(lint_ADDR_int[13]),.T1I3(lint_ADDR_int[12]),.TB1S(GND),.C1Z(NET_311),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_K6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000000000000),.B2I0(NET_142),.B2I1(GND),.B2I2(NET_141),.B2I3(NET_151),.B2Z(nx18281z1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K6_3 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_WEN_int),.T3I1(lint_ADDR_int[14]),.T3I2(lint_ADDR_int[13]),.T3I3(lint_ADDR_int[12]),.TB3S(GND),.C3Z(NET_151),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K7_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(m0_m0_dataout_int[0]),.B0I1(NET_89),.B0I2(NET_95),.B0I3(tcdm_result_p0[0]),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[12]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T0I0(m0_m0_dataout_int[0]),.T0I1(NET_89),.T0I2(NET_95),.T0I3(tcdm_result_p0[0]),.TB0S(NET_15),.C0Z(NET_113),.Q0Z(tcdm_result_p0[12]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K7_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B1I0(m0_m0_dataout_int[12]),.B1I1(NET_95),.B1I2(tcdm_result_p0[12]),.B1I3(NET_89),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[0]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p0[12]),.T1I1(NET_89),.T1I2(m0_m0_dataout_int[12]),.T1I3(NET_95),.TB1S(NET_15),.C1Z(NET_226),.Q1Z(tcdm_result_p0[0]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_K7_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B2I0(tcdm_result_p0[2]),.B2I1(NET_89),.B2I2(NET_95),.B2I3(m0_m0_dataout_int[2]),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[2]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p0[2]),.T2I1(NET_89),.T2I2(NET_95),.T2I3(m0_m0_dataout_int[2]),.TB2S(NET_15),.C2Z(NET_718),.Q2Z(tcdm_result_p0[2]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_K7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B3I0(lint_ADDR_int[2]),.B3I1(lint_ADDR_int[11]),.B3I2(apb_fsm[0]),.B3I3(lint_ADDR_int[7]),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[5]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(apb_fsm[0]),.T3I1(lint_ADDR_int[7]),.T3I2(lint_ADDR_int[2]),.T3I3(lint_ADDR_int[11]),.TB3S(lint_ADDR_int[8]),.C3Z(NET_95),.Q3Z(tcdm_result_p0[5]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q0Z(m0_m0_mode_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K8_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[6]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[12]),.T1I1(apb_fsm[0]),.T1I2(lint_ADDR_int[13]),.T1I3(GND),.C1Z(NET_41),.Q1Z(tcdm_result_p0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K8_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_89),.B2I1(NET_95),.B2I2(tcdm_result_p0[6]),.B2I3(m0_m0_dataout_int[6]),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[7]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_89),.T2I1(NET_95),.T2I2(tcdm_result_p0[6]),.T2I3(m0_m0_dataout_int[6]),.TB2S(NET_15),.C2Z(NET_636),.Q2Z(tcdm_result_p0[7]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_K8_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B3I0(tcdm_result_p0[7]),.B3I1(NET_89),.B3I2(m0_m0_dataout_int[7]),.B3I3(NET_95),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_dataout_int[7]),.T3I1(NET_95),.T3I2(tcdm_result_p0[7]),.T3I3(NET_89),.TB3S(NET_15),.C3Z(NET_470),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_K9_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_638),.B0I1(NET_639),.B0I2(NET_637),.B0I3(NET_636),.T0I0(NET_43),.T0I1(m0_coef_rdata_int[6]),.T0I2(NET_41),.T0I3(m1_coef_rdata_int[6]),.TB0S(GND),.B0Z(NET_633),.C0Z(NET_638),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K9_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_718),.T1I1(NET_719),.T1I2(NET_720),.T1I3(NET_721),.TB1S(GND),.C1Z(NET_715),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_K9_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_114),.B2I1(NET_116),.B2I2(NET_115),.B2I3(NET_113),.T2I0(NET_43),.T2I1(NET_41),.T2I2(m0_coef_rdata_int[2]),.T2I3(m1_coef_rdata_int[2]),.TB2S(GND),.B2Z(NET_105),.C2Z(NET_720),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_K9_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_43),.T3I1(m0_coef_rdata_int[0]),.T3I2(NET_41),.T3I3(m1_coef_rdata_int[0]),.TB3S(GND),.C3Z(NET_115),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K10_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_44),.T1I1(m0_oper0_rdata_int[18]),.T1I2(m1_oper1_rdata_int[18]),.T1I3(NET_117),.C1Z(NET_365),.Q1Z(m0_m1_control[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000011000000),.B2I0(NET_124),.B2I1(NET_364),.B2I2(NET_365),.B2I3(tcdm_rdata_p0_int[18]),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_124),.T2I1(NET_364),.T2I2(NET_365),.T2I3(tcdm_rdata_p0_int[18]),.TB2S(NET_366),.C2Z(NET_349),.Q2Z(m0_m0_outsel_dup_0[5]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_K10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_tc_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K11_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(m0_m0_outsel_dup_0[0]),.B0I1(tcdm_rdata_p2_int[0]),.B0I2(NET_108),.B0I3(NET_109),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p2_int[7]),.T0I1(m0_m0_control[7]),.T0I2(NET_108),.T0I3(NET_109),.TB0S(GND),.B0Z(NET_106),.C0Z(NET_468),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K11_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_8),.T1I1(GND),.T1I2(NET_38),.T1I3(lint_ADDR_int[11]),.C1Z(NET_108),.Q1Z(m0_m0_control[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K11_2 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(tcdm_rdata_p2_int[6]),.B2I1(m0_m0_tc_dup_0),.B2I2(NET_108),.B2I3(NET_109),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(NET_15),.T2I2(GND),.T2I3(NET_95),.TB2S(GND),.B2Z(NET_634),.C2Z(NET_334),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K11_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p2_int[12]),.T3I1(NET_108),.T3I2(m0_m0_mode_dup_0[0]),.T3I3(NET_109),.TB3S(GND),.C3Z(NET_224),.Q3Z(m0_m1_control[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(m0_m0_dataout_int[28]),.B0I1(NET_82),.B0I2(NET_334),.B0I3(tcdm_result_p2[28]),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(m0_m0_dataout_int[28]),.T0I1(NET_82),.T0I2(NET_334),.T0I3(tcdm_result_p2[28]),.TB0S(NET_553),.C0Z(NET_551),.Q0Z(m0_m1_control[23]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B1I0(NET_334),.B1I1(tcdm_result_p2[24]),.B1I2(m0_m0_dataout_int[24]),.B1I3(NET_82),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(m0_m0_dataout_int[24]),.T1I1(NET_82),.T1I2(NET_334),.T1I3(tcdm_result_p2[24]),.TB1S(NET_482),.C1Z(NET_480),.Q1Z(m0_m1_control[22]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_K12_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B2I0(tcdm_rdata_p2_int[22]),.B2I1(NET_109),.B2I2(m0_m1_control[22]),.B2I3(NET_112),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_112),.T2I1(NET_109),.T2I2(tcdm_rdata_p2_int[23]),.T2I3(m0_m1_control[23]),.TB2S(GND),.B2Z(NET_432),.C2Z(NET_450),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K12_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(m0_m1_control[28]),.T3I1(NET_109),.T3I2(tcdm_rdata_p2_int[28]),.T3I3(NET_112),.C3Z(NET_560),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_K13_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(NET_109),.T0I1(NET_112),.T0I2(m0_m1_control[21]),.T0I3(tcdm_rdata_p2_int[21]),.TB0S(GND),.C0Z(NET_414),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K13_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p2_int[24]),.T1I1(NET_109),.T1I2(NET_112),.T1I3(m0_m1_control[24]),.C1Z(NET_489),.Q1Z(m0_m1_control[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(tcdm_result_p3[22]),.B2I1(NET_96),.B2I2(fpgaio_out_dup_0[54]),.B2I3(NET_99),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p3[22]),.T2I1(NET_96),.T2I2(fpgaio_out_dup_0[54]),.T2I3(NET_99),.TB2S(NET_429),.C2Z(NET_426),.Q2Z(m0_coef_wmode_dup_0[0]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_K13_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(NET_109),.T3I1(tcdm_rdata_p2_int[2]),.T3I2(NET_108),.T3I3(m0_m0_outsel_dup_0[2]),.TB3S(GND),.C3Z(NET_716),.Q3Z(m0_m1_control[21]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K14_0 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_326),.B0I1(NET_328),.B0I2(NET_327),.B0I3(NET_329),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.T0I0(lint_ADDR_int[14]),.T0I1(apb_fsm[0]),.T0I2(GND),.T0I3(lint_ADDR_int[12]),.TB0S(GND),.B0Z(NET_313),.C0Z(NET_44),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K14_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.T1I0(tcdm_rdata_p2_int[16]),.T1I1(m0_m0_rnd_dup_0),.T1I2(NET_6),.T1I3(NET_36),.C1Z(NET_329),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K14_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_156),.B2I1(NET_729),.B2I2(NET_164),.B2I3(NET_161),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.T2I0(NET_156),.T2I1(NET_729),.T2I2(NET_164),.T2I3(NET_161),.TB2S(NET_170),.Q2Z(lint_RDATA_dup_0[9]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_K14_3 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.T3I0(GND),.T3I1(NET_8),.T3I2(GND),.T3I3(NET_38),.TB3S(GND),.C3Z(NET_36),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_K15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000010000000),.B0I0(lint_WEN_int),.B0I1(lint_ADDR_int[14]),.B0I2(lint_ADDR_int[13]),.B0I3(lint_ADDR_int[12]),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.B0Z(NET_140),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K15_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[5]),.T1I1(lint_ADDR_int[6]),.T1I2(NET_134),.T1I3(NET_146),.TB1S(GND),.C1Z(nx19726z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_K15_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[11]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_598),.T2I1(NET_600),.T2I2(NET_599),.T2I3(NET_601),.TB2S(GND),.C2Z(NET_586),.Q2Z(tcdm_result_p0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_K15_3 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(lint_WEN_int),.T3I1(lint_ADDR_int[14]),.T3I2(lint_ADDR_int[13]),.T3I3(lint_ADDR_int[12]),.TB3S(GND),.C3Z(NET_645),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_K16_0 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0001000000000000),.B0I0(GND),.B0I1(GND),.B0I2(NET_8),.B0I3(NET_7),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(NET_69),.T0I2(lint_ADDR_int[4]),.T0I3(NET_70),.TB0S(GND),.B0Z(NET_6),.C0Z(NET_67),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K16_1 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[7]),.T1I1(lint_ADDR_int[2]),.T1I2(NET_15),.T1I3(NET_19),.TB1S(GND),.C1Z(NET_59),.Q1Z(m0_m0_outsel_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_K16_2 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0001000000000000),.B2I0(GND),.B2I1(GND),.B2I2(NET_7),.B2I3(NET_95),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[6]),.T2I1(NET_11),.T2I2(NET_8),.T2I3(lint_ADDR_int[5]),.TB2S(GND),.B2Z(NET_94),.C2Z(NET_61),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K16_3 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(lint_ADDR_int[11]),.T3I2(NET_11),.T3I3(lint_ADDR_int[7]),.TB3S(GND),.C3Z(NET_148),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_K17_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_686),.B0I1(NET_688),.B0I2(NET_689),.B0I3(NET_687),.T0I0(NET_160),.T0I1(NET_157),.T0I2(NET_159),.T0I3(NET_158),.TB0S(GND),.B0Z(NET_690),.C0Z(NET_161),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K17_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(GND),.T1I1(lint_ADDR_int[4]),.T1I2(GND),.T1I3(lint_ADDR_int[3]),.TB1S(GND),.C1Z(NET_11),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_K17_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.T2I0(fpgaio_out_dup_0[35]),.T2I1(NET_6),.T2I2(tcdm_rdata_p2_int[3]),.T2I3(NET_5),.TB2S(GND),.C2Z(NET_688),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_K17_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_12),.T3I1(NET_13),.T3I2(tcdm_result_p0[3]),.T3I3(fpgaio_out_dup_0[67]),.TB3S(GND),.C3Z(NET_689),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K18_0 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_13),.B0I1(tcdm_result_p0[5]),.B0I2(fpgaio_out_dup_0[69]),.B0I3(NET_12),.T0I0(NET_11),.T0I1(lint_ADDR_int[6]),.T0I2(lint_ADDR_int[5]),.T0I3(NET_10),.TB0S(GND),.B0Z(NET_650),.C0Z(NET_17),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K18_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_153),.T1I1(NET_155),.T1I2(NET_154),.T1I3(NET_152),.C1Z(NET_156),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K18_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_13),.B2I1(tcdm_result_p0[9]),.B2I2(NET_12),.B2I3(fpgaio_out_dup_0[73]),.T2I0(NET_5),.T2I1(fpgaio_out_dup_0[40]),.T2I2(NET_6),.T2I3(tcdm_rdata_p2_int[8]),.TB2S(GND),.B2Z(NET_155),.C2Z(NET_275),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_K18_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_5),.T3I1(fpgaio_out_dup_0[41]),.T3I2(NET_6),.T3I3(tcdm_rdata_p2_int[9]),.TB3S(GND),.C3Z(NET_154),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K19_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B0I0(m1_m0_dataout_int[3]),.B0I1(m1_ram_control[3]),.B0I2(NET_17_CAND2_BLSTR_11_tpGCLKBUF),.B0I3(NET_18_CAND4_BLSTR_11_tpGCLKBUF),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T0I0(NET_61),.T0I1(m1_m0_dataout_int[20]),.T0I2(m0_ram_control[20]),.T0I3(NET_18_CAND4_BLSTR_11_tpGCLKBUF),.TB0S(GND),.B0Z(NET_687),.C0Z(NET_400),.Q0Z(m0_ram_control[31]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q1Z(m0_ram_control[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K19_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000001000),.B2I0(NET_19),.B2I1(NET_7),.B2I2(lint_ADDR_int[2]),.B2I3(lint_ADDR_int[7]),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx49871z1_CAND3_BLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_61),.T2I1(m1_m0_dataout_int[31]),.T2I2(NET_18_CAND4_BLSTR_11_tpGCLKBUF),.T2I3(m0_ram_control[31]),.TB2S(GND),.B2Z(NET_18),.C2Z(NET_617),.Q2Z(m1_ram_control[3]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_K19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdsel_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K20_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T0I0(m1_m0_dataout_int[27]),.T0I1(NET_18_CAND4_BLSTR_11_tpGCLKBUF),.T0I2(m0_ram_control[27]),.T0I3(NET_61),.TB0S(GND),.C0Z(NET_546),.Q0Z(m0_ram_control[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q1Z(m0_ram_control[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K20_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(m0_ram_control[30]),.T3I1(m1_m0_dataout_int[30]),.T3I2(NET_18_CAND4_BLSTR_11_tpGCLKBUF),.T3I3(NET_61),.TB3S(GND),.C3Z(NET_599),.Q3Z(m0_oper1_rmode_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_rmode_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K21_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_18_CAND4_BLSTR_11_tpGCLKBUF),.T1I1(m1_m0_dataout_int[9]),.T1I2(m1_ram_control[9]),.T1I3(NET_17_CAND2_BLSTR_11_tpGCLKBUF),.TB1S(GND),.C1Z(NET_153),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_K21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_m0_dataout_int[1]),.B2I1(m1_ram_control[1]),.B2I2(NET_18_CAND4_BLSTR_11_tpGCLKBUF),.B2I3(NET_17_CAND2_BLSTR_11_tpGCLKBUF),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx49871z1_CAND3_BLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.B2Z(NET_1),.Q2Z(m1_ram_control[1]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx49871z1_CAND3_BLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q3Z(m1_ram_control[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m1_m1_dataout_int[9]),.B0I1(NET_33),.B0I2(m1_m0_control[9]),.B0I3(NET_32),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B0Z(NET_160),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K26_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_253),.T1I1(NET_143),.T1I2(lint_ADDR_int[13]),.T1I3(NET_65),.TB1S(GND),.C1Z(nx30664z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_K26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_control[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_65),.B2I1(lint_ADDR_int[13]),.B2I2(GND),.B2I3(NET_171),.B2Z(nx33579z1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K29_0 (.tFragBitInfo(16'b0000000000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(apb_fsm[0]),.T0I1(lint_ADDR_int[12]),.T0I2(lint_ADDR_int[13]),.T0I3(GND),.TB0S(GND),.C0Z(NET_45),.Q0Z(m1_coef_wdata_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_mode_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K30_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_32),.T1I1(NET_33),.T1I2(m1_m1_dataout_int[13]),.T1I3(m1_m0_mode_dup_0[1]),.C1Z(NET_242),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_reset_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_oper1_rdata_int[0]),.B2I1(NET_45_CAND5_BLSBR_11_tpGCLKBUF),.B2I2(NET_44_CAND4_BLSBR_11_tpGCLKBUF),.B2I3(m1_oper0_rdata_int[0]),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B2Z(NET_116),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K31_3 (.tFragBitInfo(16'b1111001111110011),.bFragBitInfo(16'b1010100011111101),.B3I0(apb_fsm[0]),.B3I1(lint_ADDR_int[12]),.B3I2(lint_ADDR_int[13]),.B3I3(lint_ADDR_int[11]),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[13]),.T3I1(lint_ADDR_int[11]),.T3I2(apb_fsm[0]),.T3I3(lint_ADDR_int[12]),.TB3S(m1_oper0_rdata_int[16]),.C3Z(NET_742),.Q3Z(m1_coef_wdata_dup_0[31]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K32_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_45_CAND5_BLSBR_11_tpGCLKBUF),.B0I1(m1_oper1_rdata_int[2]),.B0I2(NET_44_CAND4_BLSBR_11_tpGCLKBUF),.B0I3(m1_oper0_rdata_int[2]),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(m1_coef_rdata_int[26]),.T0I1(m1_oper0_rdata_int[26]),.T0I2(NET_43_CAND3_BLSBR_11_tpGCLKBUF),.T0I3(NET_45_CAND5_BLSBR_11_tpGCLKBUF),.TB0S(GND),.B0Z(NET_721),.C0Z(NET_528),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K32_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[21]),.Q1EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(m1_coef_rdata_int[17]),.T1I1(m1_oper0_rdata_int[17]),.T1I2(NET_43_CAND3_BLSBR_11_tpGCLKBUF),.T1I3(NET_45_CAND5_BLSBR_11_tpGCLKBUF),.TB1S(GND),.C1Z(NET_346),.Q1Z(m1_coef_wdata_dup_0[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_K32_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_45_CAND5_BLSBR_11_tpGCLKBUF),.T2I1(NET_43_CAND3_BLSBR_11_tpGCLKBUF),.T2I2(m1_coef_rdata_int[23]),.T2I3(m1_oper0_rdata_int[23]),.TB2S(GND),.C2Z(NET_454),.Q2Z(m1_coef_wdata_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_K32_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(m1_oper0_rdata_int[6]),.T3I1(NET_45_CAND5_BLSBR_11_tpGCLKBUF),.T3I2(m1_oper1_rdata_int[6]),.T3I3(NET_44_CAND4_BLSBR_11_tpGCLKBUF),.TB3S(GND),.C3Z(NET_639),.Q3Z(m1_coef_wdata_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[21]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L6_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_141),.T1I1(GND),.T1I2(NET_311),.T1I3(NET_142),.C1Z(nx32231z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_L6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L8_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[14]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.T0I0(NET_62),.T0I1(NET_63),.T0I2(tcdm_rdata_p0_int[10]),.T0I3(m0_m1_control[10]),.TB0S(GND),.C0Z(NET_190),.Q0Z(tcdm_result_p0[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[9]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_control[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L8_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_62),.T3I1(NET_63),.T3I2(m0_m1_control[9]),.T3I3(tcdm_rdata_p0_int[9]),.TB3S(GND),.C3Z(NET_167),.Q3Z(m0_m1_control[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L9_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(NET_62),.T0I1(tcdm_rdata_p0_int[8]),.T0I2(NET_63),.T0I3(m0_m1_control[8]),.TB0S(GND),.C0Z(NET_288),.Q0Z(m0_m1_control[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.Q2Z(m0_m0_reset_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[8]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L10_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000100000),.B0I0(NET_38),.B0I1(lint_ADDR_int[11]),.B0I2(NET_10),.B0I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(NET_117),.T0I1(m0_oper0_rdata_int[22]),.T0I2(m1_oper1_rdata_int[22]),.T0I3(NET_44),.TB0S(GND),.B0Z(NET_112),.C0Z(NET_437),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L10_1 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[9]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_38),.T1I1(GND),.T1I2(GND),.T1I3(NET_10),.TB1S(GND),.C1Z(NET_63),.Q1Z(tcdm_result_p0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_L10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000100),.B2I0(lint_ADDR_int[5]),.B2I1(lint_ADDR_int[4]),.B2I2(lint_ADDR_int[3]),.B2I3(lint_ADDR_int[6]),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.B2Z(NET_38),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000011000000),.B3I0(tcdm_rdata_p0_int[22]),.B3I1(NET_437),.B3I2(NET_436),.B3I3(NET_124),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_436),.T3I1(NET_124),.T3I2(tcdm_rdata_p0_int[22]),.T3I3(NET_437),.TB3S(NET_438),.C3Z(NET_421),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_L11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_82),.B0I1(m0_m0_dataout_int[23]),.B0I2(NET_334),.B0I3(tcdm_result_p2[23]),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[10]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(NET_82),.T0I1(m0_m0_dataout_int[23]),.T0I2(NET_334),.T0I3(tcdm_result_p2[23]),.TB0S(NET_443),.C0Z(NET_441),.Q0Z(tcdm_result_p0[10]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B1I0(tcdm_result_p2[19]),.B1I1(m0_m0_dataout_int[19]),.B1I2(NET_82),.B1I3(NET_334),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[23]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_82),.T1I1(NET_334),.T1I2(tcdm_result_p2[19]),.T1I3(m0_m0_dataout_int[19]),.TB1S(NET_372),.C1Z(NET_370),.Q1Z(tcdm_result_p2[23]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_L11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_82),.B2I1(m0_m0_dataout_int[26]),.B2I2(NET_334),.B2I3(tcdm_result_p2[26]),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T2I0(NET_82),.T2I1(m0_m0_dataout_int[26]),.T2I2(NET_334),.T2I3(tcdm_result_p2[26]),.TB2S(NET_517),.C2Z(NET_515),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_L11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B3I0(NET_334),.B3I1(m0_m0_dataout_int[29]),.B3I2(NET_82),.B3I3(tcdm_result_p2[29]),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[19]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_82),.T3I1(tcdm_result_p2[29]),.T3I2(NET_334),.T3I3(m0_m0_dataout_int[29]),.TB3S(NET_571),.C3Z(NET_569),.Q3Z(tcdm_result_p2[19]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_82),.B0I1(m0_m0_dataout_int[18]),.B0I2(tcdm_result_p2[18]),.B0I3(NET_334),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[24]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(NET_82),.T0I1(m0_m0_dataout_int[18]),.T0I2(tcdm_result_p2[18]),.T0I3(NET_334),.TB0S(NET_353),.C0Z(NET_351),.Q0Z(tcdm_result_p2[24]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(m0_m0_dataout_int[22]),.B1I1(NET_334),.B1I2(NET_82),.B1I3(tcdm_result_p2[22]),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[28]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_82),.T1I1(tcdm_result_p2[22]),.T1I2(m0_m0_dataout_int[22]),.T1I3(NET_334),.TB1S(NET_425),.C1Z(NET_423),.Q1Z(tcdm_result_p2[28]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_L12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_82),.B2I1(tcdm_result_p2[17]),.B2I2(NET_334),.B2I3(m0_m0_dataout_int[17]),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[22]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T2I0(NET_82),.T2I1(tcdm_result_p2[17]),.T2I2(NET_334),.T2I3(m0_m0_dataout_int[17]),.TB2S(NET_335),.C2Z(NET_332),.Q2Z(tcdm_result_p2[22]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_L12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(tcdm_result_p2[21]),.B3I1(NET_334),.B3I2(NET_82),.B3I3(m0_m0_dataout_int[21]),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[21]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_82),.T3I1(m0_m0_dataout_int[21]),.T3I2(tcdm_result_p2[21]),.T3I3(NET_334),.TB3S(NET_407),.C3Z(NET_405),.Q3Z(tcdm_result_p2[21]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L14_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_313),.B0I1(NET_312),.B0I2(NET_314),.B0I3(NET_315),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T0I0(NET_313),.T0I1(NET_312),.T0I2(NET_314),.T0I3(NET_315),.TB0S(NET_316),.Q0Z(lint_RDATA_dup_0[16]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L14_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T1I0(tcdm_rdata_p2_int[31]),.T1I1(NET_36),.T1I2(NET_6),.T1I3(m0_m0_reset_dup_0),.TB1S(GND),.C1Z(NET_619),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(tcdm_result_p3[29]),.B2I1(fpgaio_out_dup_0[61]),.B2I2(NET_96),.B2I3(NET_99),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T2I0(tcdm_result_p3[29]),.T2I1(fpgaio_out_dup_0[61]),.T2I2(NET_96),.T2I3(NET_99),.TB2S(NET_575),.C2Z(NET_572),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_L14_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T3I0(NET_617),.T3I1(NET_616),.T3I2(NET_619),.T3I3(NET_618),.C3Z(NET_604),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L15_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_588),.B0I1(NET_587),.B0I2(NET_586),.B0I3(NET_585),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T0I0(NET_588),.T0I1(NET_587),.T0I2(NET_586),.T0I3(NET_585),.TB0S(NET_589),.Q0Z(lint_RDATA_dup_0[30]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L15_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T1I0(NET_545),.T1I1(NET_547),.T1I2(NET_548),.T1I3(NET_546),.TB1S(GND),.C1Z(NET_533),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L15_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000010000000),.B2I0(NET_140),.B2I1(NET_141),.B2I2(NET_142),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T2I0(NET_141),.T2I1(NET_645),.T2I2(NET_142),.T2I3(GND),.TB2S(GND),.B2Z(nx14650z1),.C2Z(nx53672z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_L15_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T3I0(NET_512),.T3I1(NET_510),.T3I2(NET_511),.T3I3(NET_509),.TB3S(GND),.C3Z(NET_497),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_L16_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_36),.B0I1(NET_6),.B0I2(m0_m0_control[20]),.B0I3(tcdm_rdata_p2_int[20]),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(m0_m0_control[27]),.T0I1(NET_6),.T0I2(tcdm_rdata_p2_int[27]),.T0I3(NET_36),.TB0S(GND),.B0Z(NET_402),.C0Z(NET_548),.Q0Z(m0_m0_control[25]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L16_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_401),.T1I1(NET_399),.T1I2(NET_402),.T1I3(NET_400),.C1Z(NET_387),.Q1Z(m0_m0_control[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_L16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_36),.B2I1(NET_6),.B2I2(m0_m0_control[30]),.B2I3(tcdm_rdata_p2_int[30]),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.B2Z(NET_601),.Q2Z(m0_m0_control[27]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L16_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_36),.T3I1(NET_6),.T3I2(tcdm_rdata_p2_int[25]),.T3I3(m0_m0_control[25]),.TB3S(GND),.C3Z(NET_512),.Q3Z(m0_m0_control[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_clr_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_control[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_590),.B2I1(NET_591),.B2I2(NET_593),.B2I3(NET_592),.CD2S(VCC),.Q2DI(lint_WDATA_int[30]),.Q2EN(nx49871z1_CAND3_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B2Z(NET_587),.Q2Z(m1_ram_control[30]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L18_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.B3I0(m1_m1_control[30]),.B3I1(NET_17_CAND2_BLSTR_12_tpGCLKBUF),.B3I2(NET_28_CAND5_BLSTR_12_tpGCLKBUF),.B3I3(m1_ram_control[30]),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_28_CAND5_BLSTR_12_tpGCLKBUF),.T3I1(m1_ram_control[30]),.T3I2(m1_m1_control[30]),.T3I3(NET_17_CAND2_BLSTR_12_tpGCLKBUF),.TB3S(NET_594),.C3Z(NET_592),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_L19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L19_1 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[7]),.T1I1(NET_19),.T1I2(lint_ADDR_int[2]),.T1I3(NET_7),.C1Z(NET_33),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_L19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L19_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_539),.T3I1(NET_538),.T3I2(NET_540),.T3I3(NET_537),.C3Z(NET_534),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m1_m1_dataout_int[27]),.B0I1(NET_33),.B0I2(NET_32),.B0I3(m1_m0_control[27]),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B0Z(NET_538),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q3Z(m1_m0_control[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m1_m0_control[11]),.B0I1(NET_32),.B0I2(m1_m1_dataout_int[11]),.B0I3(NET_33),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.B0Z(NET_202),.Q0Z(m1_m0_control[11]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[22]),.Q0EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[25]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L32_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(m1_coef_rdata_int[10]),.T0I1(NET_43_CAND3_BLSBR_12_tpGCLKBUF),.T0I2(NET_44_CAND4_BLSBR_12_tpGCLKBUF),.T0I3(m1_oper1_rdata_int[10]),.TB0S(GND),.C0Z(NET_185),.Q0Z(m1_coef_wdata_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L32_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_44_CAND4_BLSBR_12_tpGCLKBUF),.T1I1(NET_43_CAND3_BLSBR_12_tpGCLKBUF),.T1I2(m1_coef_rdata_int[13]),.T1I3(m1_oper1_rdata_int[13]),.TB1S(GND),.C1Z(NET_244),.Q1Z(m1_coef_wdata_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_L32_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_rdata_int[14]),.T2I1(NET_43_CAND3_BLSBR_12_tpGCLKBUF),.T2I2(m1_coef_rdata_int[14]),.T2I3(NET_44_CAND4_BLSBR_12_tpGCLKBUF),.TB2S(GND),.C2Z(NET_264),.Q2Z(m1_coef_wdata_dup_0[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_L32_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[20]),.Q3EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(m1_oper1_rdata_int[11]),.T3I1(m1_coef_rdata_int[11]),.T3I2(NET_44_CAND4_BLSBR_12_tpGCLKBUF),.T3I3(NET_43_CAND3_BLSBR_12_tpGCLKBUF),.TB3S(GND),.C3Z(NET_204),.Q3Z(m1_coef_wdata_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M1_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[4]),.Q0EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(m0_coef_rdata_int[22]),.T0I1(NET_41_CAND4_TLSTR_13_tpGCLKBUF),.T0I2(m0_oper1_rdata_int[22]),.T0I3(NET_46_CAND3_TLSTR_13_tpGCLKBUF),.TB0S(GND),.C0Z(NET_438),.Q0Z(m0_coef_waddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[9]),.Q1EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_waddr_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[10]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_waddr_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[5]),.Q1EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_waddr_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[11]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_waddr_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_outsel_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M7_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_62),.T3I1(NET_63),.T3I2(tcdm_rdata_p0_int[14]),.T3I3(m0_m1_osel_dup_0),.TB3S(GND),.C3Z(NET_269),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_M8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(lint_ADDR_int[11]),.B0I1(apb_fsm[0]),.B0I2(lint_ADDR_int[8]),.B0I3(lint_ADDR_int[2]),.CD0S(VCC),.Q0DI(lint_WDATA_int[17]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[11]),.T0I1(apb_fsm[0]),.T0I2(lint_ADDR_int[8]),.T0I3(lint_ADDR_int[2]),.TB0S(lint_ADDR_int[7]),.C0Z(NET_89),.Q0Z(m0_m1_clr_dup_0),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_m0_outsel_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[4]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[13]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M10_0 (.tFragBitInfo(16'b1010000000000000),.bFragBitInfo(16'b0010000000000000),.B0I0(NET_397),.B0I1(m0_oper0_rdata_int[20]),.B0I2(NET_745),.B0I3(NET_398),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_397),.T0I1(m0_oper0_rdata_int[20]),.T0I2(NET_745),.T0I3(NET_398),.TB0S(NET_117),.C0Z(NET_389),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_control[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M10_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_44),.B2I1(NET_117),.B2I2(m1_oper1_rdata_int[21]),.B2I3(m0_oper0_rdata_int[21]),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_63),.T2I1(NET_62),.T2I2(tcdm_rdata_p0_int[11]),.T2I3(m0_m1_control[11]),.TB2S(GND),.B2Z(NET_419),.C2Z(NET_209),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_M10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100110000000000),.B3I0(tcdm_rdata_p0_int[21]),.B3I1(NET_418),.B3I2(NET_124),.B3I3(NET_419),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_124),.T3I1(NET_419),.T3I2(tcdm_rdata_p0_int[21]),.T3I3(NET_418),.TB3S(NET_420),.C3Z(NET_403),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_M11_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000010000000000),.B0I0(GND),.B0I1(NET_8),.B0I2(GND),.B0I3(NET_125_CAND4_TLSBR_13_tpGCLKBUF),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_109),.T0I1(tcdm_rdata_p2_int[29]),.T0I2(NET_112),.T0I3(m0_m1_control[29]),.TB0S(GND),.B0Z(NET_124),.C0Z(NET_578),.Q0Z(m0_m1_control[29]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M11_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[26]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(m0_oper0_rdata_int[19]),.T1I1(m1_oper1_rdata_int[19]),.T1I2(NET_117),.T1I3(NET_44),.TB1S(GND),.C1Z(NET_384),.Q1Z(tcdm_result_p2[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[29]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p2[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000010100000),.B3I0(NET_384),.B3I1(tcdm_rdata_p0_int[19]),.B3I2(NET_383),.B3I3(NET_124),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_383),.T3I1(NET_124),.T3I2(NET_384),.T3I3(tcdm_rdata_p0_int[19]),.TB3S(NET_385),.C3Z(NET_368),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_M12_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B0I0(tcdm_rdata_p3_int[18]),.B0I1(NET_110_CAND3_TLSBR_13_tpGCLKBUF),.B0I2(tcdm_rdata_p1_int[18]),.B0I3(NET_125_CAND4_TLSBR_13_tpGCLKBUF),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[18]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p3_int[18]),.T0I1(NET_110_CAND3_TLSBR_13_tpGCLKBUF),.T0I2(tcdm_rdata_p1_int[18]),.T0I3(NET_125_CAND4_TLSBR_13_tpGCLKBUF),.TB0S(NET_10),.C0Z(NET_363),.Q0Z(tcdm_result_p2[18]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M12_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[17]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_66),.T1I1(NET_145),.T1I2(GND),.T1I3(NET_67),.TB1S(GND),.C1Z(nx40728z1),.Q1Z(tcdm_result_p2[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m0_m1_clr_dup_0),.B2I1(tcdm_rdata_p2_int[17]),.B2I2(NET_112),.B2I3(NET_109),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B2Z(NET_342),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M12_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(m0_m1_sat_dup_0),.T3I1(tcdm_rdata_p2_int[18]),.T3I2(NET_112),.T3I3(NET_109),.C3Z(NET_360),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_99),.B0I1(fpgaio_out_dup_0[55]),.B0I2(NET_96),.B0I3(tcdm_result_p3[23]),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_99),.T0I1(fpgaio_out_dup_0[55]),.T0I2(NET_96),.T0I3(tcdm_result_p3[23]),.TB0S(NET_447),.C0Z(NET_444),.Q0Z(m0_m1_control[19]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M13_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_112),.T1I1(NET_109),.T1I2(tcdm_rdata_p2_int[19]),.T1I3(m0_m1_control[19]),.C1Z(NET_379),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_M13_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000001000000000),.B2I0(NET_110_CAND3_TLSBR_13_tpGCLKBUF),.B2I1(GND),.B2I2(GND),.B2I3(NET_8),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p2_int[26]),.T2I1(NET_109),.T2I2(m0_m1_control[26]),.T2I3(NET_112),.TB2S(GND),.B2Z(NET_109),.C2Z(NET_524),.Q2Z(m0_m1_control[26]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_M13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B3I0(NET_96),.B3I1(tcdm_result_p3[17]),.B3I2(NET_99),.B3I3(fpgaio_out_dup_0[49]),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_99),.T3I1(fpgaio_out_dup_0[49]),.T3I2(NET_96),.T3I3(tcdm_result_p3[17]),.TB3S(NET_339),.C3Z(NET_336),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_M14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(fpgaio_out_dup_0[60]),.B0I1(NET_96),.B0I2(tcdm_result_p3[28]),.B0I3(NET_99),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.T0I0(fpgaio_out_dup_0[60]),.T0I1(NET_96),.T0I2(tcdm_result_p3[28]),.T0I3(NET_99),.TB0S(NET_557),.C0Z(NET_554),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M14_1 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.T1I0(NET_8),.T1I1(NET_15),.T1I2(GND),.T1I3(GND),.TB1S(GND),.C1Z(NET_62),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_M14_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_606),.B2I1(NET_604),.B2I2(NET_603),.B2I3(NET_605),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.T2I0(NET_606),.T2I1(NET_604),.T2I2(NET_603),.T2I3(NET_605),.TB2S(NET_607),.Q2Z(lint_RDATA_dup_0[31]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_M14_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_386),.B3I1(NET_387),.B3I2(NET_388),.B3I3(NET_389),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.T3I0(NET_388),.T3I1(NET_389),.T3I2(NET_386),.T3I3(NET_387),.TB3S(NET_390),.Q3Z(lint_RDATA_dup_0[20]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_M15_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_499),.B0I1(NET_497),.B0I2(NET_496),.B0I3(NET_498),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.T0I0(NET_499),.T0I1(NET_497),.T0I2(NET_496),.T0I3(NET_498),.TB0S(NET_500),.Q0Z(lint_RDATA_dup_0[25]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M15_1 (.tFragBitInfo(16'b1101110011011100),.bFragBitInfo(16'b1111111100001110),.B1I0(NET_147),.B1I1(NET_755),.B1I2(nx7012z3),.B1I3(NET_621),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.T1I0(nx7012z3),.T1I1(NET_621),.T1I2(NET_147),.T1I3(NET_755),.TB1S(NET_69),.C1Z(nx49808z64),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_M15_2 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b0000001000000000),.B2I0(NET_148),.B2I1(GND),.B2I2(GND),.B2I3(NET_69),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.T2I0(NET_148),.T2I1(NET_65),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(NET_146),.C2Z(NET_174),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_M15_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_534),.B3I1(NET_532),.B3I2(NET_535),.B3I3(NET_533),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.T3I0(NET_535),.T3I1(NET_533),.T3I2(NET_534),.T3I3(NET_532),.TB3S(NET_536),.Q3Z(lint_RDATA_dup_0[27]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_M16_0 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_65),.B0I1(NET_68),.B0I2(NET_66),.B0I3(NET_67),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(lint_ADDR_int[2]),.T0I2(lint_ADDR_int[11]),.T0I3(NET_75),.TB0S(GND),.B0Z(nx10775z1),.C0Z(NET_76),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M16_1 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[3]),.T1I1(lint_ADDR_int[11]),.T1I2(GND),.T1I3(NET_75),.TB1S(GND),.C1Z(NET_70),.Q1Z(m0_m0_outsel_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M16_2 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_76),.T2I1(NET_69),.T2I2(GND),.T2I3(GND),.TB2S(GND),.C2Z(NET_68),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_M16_3 (.tFragBitInfo(16'b1111111111111011),.bFragBitInfo(16'b1111111111111111),.B3I0(NET_70),.B3I1(NET_62),.B3I2(NET_76),.B3I3(NET_754),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_76),.T3I1(NET_754),.T3I2(NET_70),.T3I3(NET_62),.TB3S(NET_148),.C3Z(NET_755),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_M17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_68),.B0I1(NET_66),.B0I2(lint_ADDR_int[3]),.B0I3(NET_65),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_68),.T0I1(NET_66),.T0I2(lint_ADDR_int[3]),.T0I3(NET_65),.TB0S(lint_ADDR_int[4]),.C0Z(nx28356z1),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_m1_mode_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M18_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.B0I0(NET_28_CAND5_BLSTR_13_tpGCLKBUF),.B0I1(m1_ram_control[20]),.B0I2(NET_17_CAND2_BLSTR_13_tpGCLKBUF),.B0I3(m1_m1_control[20]),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx49871z1_CAND3_BLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_28_CAND5_BLSTR_13_tpGCLKBUF),.T0I1(m1_ram_control[20]),.T0I2(NET_17_CAND2_BLSTR_13_tpGCLKBUF),.T0I3(m1_m1_control[20]),.TB0S(NET_395),.C0Z(NET_393),.Q0Z(m1_ram_control[20]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M18_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_504),.T1I1(NET_503),.T1I2(NET_502),.T1I3(NET_501),.C1Z(NET_498),.Q1Z(m1_m1_control[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_M18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_393),.B0I1(NET_392),.B0I2(NET_391),.B0I3(NET_394),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B0Z(NET_388),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M19_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.B2I0(NET_17_CAND2_BLSTR_13_tpGCLKBUF),.B2I1(m1_ram_control[27]),.B2I2(NET_28_CAND5_BLSTR_13_tpGCLKBUF),.B2I3(m1_m1_control[27]),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx49871z1_CAND3_BLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_17_CAND2_BLSTR_13_tpGCLKBUF),.T2I1(m1_ram_control[27]),.T2I2(m1_m1_control[27]),.T2I3(NET_28_CAND5_BLSTR_13_tpGCLKBUF),.TB2S(NET_541),.C2Z(NET_539),.Q2Z(m1_ram_control[27]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_M19_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_609),.T3I1(NET_611),.T3I2(NET_608),.T3I3(NET_610),.TB3S(GND),.C3Z(NET_605),.Q3Z(m1_m1_control[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_control[25]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M20_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_dataout_int[25]),.T1I1(NET_33),.T1I2(NET_32),.T1I3(m1_m0_control[25]),.C1Z(NET_502),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_M20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_control[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M21_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(m1_m1_dataout_int[20]),.T3I1(m1_m0_control[20]),.T3I2(NET_32),.T3I3(NET_33),.C3Z(NET_392),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(m1_m1_dataout_int[10]),.B0I1(NET_32),.B0I2(NET_33),.B0I3(m1_m0_control[10]),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B0Z(NET_183),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_control[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_control[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_m0_control[30]),.B2I1(NET_33),.B2I2(NET_32),.B2I3(m1_m1_dataout_int[30]),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B2Z(NET_591),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M30_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_reset_dup_0),.T3I1(NET_32),.T3I2(NET_33),.T3I3(m1_m1_dataout_int[31]),.TB3S(GND),.C3Z(NET_609),.Q3Z(m1_coef_wdata_dup_0[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[11]),.Q1EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_waddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[4]),.Q0EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_waddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M32_1 (.tFragBitInfo(16'b0100010011001100),.bFragBitInfo(16'b0001010100000000),.B1I0(m1_oper1_rdata_int[20]),.B1I1(m1_coef_rdata_int[20]),.B1I2(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.B1I3(NET_744),.CD1S(VCC),.Q1DI(lint_ADDR_int[0]),.Q1EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.T1I1(NET_744),.T1I2(m1_oper1_rdata_int[20]),.T1I3(m1_coef_rdata_int[20]),.TB1S(NET_44_CAND4_BLSBR_13_tpGCLKBUF),.C1Z(NET_745),.Q1Z(m1_coef_waddr_dup_0[0]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_44_CAND4_BLSBR_13_tpGCLKBUF),.B2I1(m1_oper1_rdata_int[9]),.B2I2(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.B2I3(m1_coef_rdata_int[9]),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B2Z(NET_162),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_waddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N1_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[0]),.Q0EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.T0I0(m0_oper1_rdata_int[28]),.T0I1(NET_46_CAND3_TLSTR_14_tpGCLKBUF),.T0I2(NET_41_CAND4_TLSTR_14_tpGCLKBUF),.T0I3(m0_coef_rdata_int[28]),.TB0S(GND),.C0Z(NET_566),.Q0Z(m0_coef_waddr_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N1_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[1]),.Q1EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_46_CAND3_TLSTR_14_tpGCLKBUF),.T1I1(m0_oper1_rdata_int[16]),.T1I2(NET_41_CAND4_TLSTR_14_tpGCLKBUF),.T1I3(m0_coef_rdata_int[16]),.TB1S(GND),.C1Z(NET_325),.Q1Z(m0_coef_waddr_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[10]),.Q2EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_raddr_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[7]),.Q3EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_waddr_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[2]),.Q0EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_waddr_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(NET_762),.Q1EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_we_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[6]),.Q2EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_waddr_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[9]),.Q3EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_raddr_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[8]),.Q0EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_raddr_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[8]),.Q1EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_waddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[3]),.Q2EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_waddr_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[11]),.Q3EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_raddr_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N4_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_65),.T1I1(NET_149),.T1I2(lint_ADDR_int[13]),.T1I3(GND),.TB1S(GND),.C1Z(nx25587z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_N4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_osel_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N7_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.T0I0(m0_m1_mode_dup_0[1]),.T0I1(NET_62),.T0I2(tcdm_rdata_p0_int[13]),.T0I3(NET_63),.TB0S(GND),.C0Z(NET_249),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_mode_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(m0_m1_outsel_dup_0[5]),.B2I1(NET_62),.B2I2(tcdm_rdata_p0_int[5]),.B2I3(NET_63),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B2Z(NET_662),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[15]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.Q0Z(m0_m1_outsel_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[1]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N10_0 (.tFragBitInfo(16'b1010000000000000),.bFragBitInfo(16'b0010000000000000),.B0I0(NET_747),.B0I1(m0_oper0_rdata_int[25]),.B0I2(NET_507),.B0I3(NET_508),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_747),.T0I1(m0_oper0_rdata_int[25]),.T0I2(NET_507),.T0I3(NET_508),.TB0S(NET_117),.C0Z(NET_499),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N10_1 (.tFragBitInfo(16'b1000100000000000),.bFragBitInfo(16'b0100000000000000),.B1I0(m0_oper0_rdata_int[16]),.B1I1(NET_325),.B1I2(NET_743),.B1I3(NET_324),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[22]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_743),.T1I1(NET_324),.T1I2(m0_oper0_rdata_int[16]),.T1I3(NET_325),.TB1S(NET_117),.C1Z(NET_315),.Q1Z(tcdm_result_p0[22]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[18]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p0[18]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N10_3 (.tFragBitInfo(16'b1000000010000000),.bFragBitInfo(16'b0010000000000000),.B3I0(NET_749),.B3I1(m0_oper0_rdata_int[27]),.B3I2(NET_543),.B3I3(NET_544),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(NET_543),.T3I1(NET_544),.T3I2(NET_749),.T3I3(m0_oper0_rdata_int[27]),.TB3S(NET_117),.C3Z(NET_535),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_N11_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_44),.B0I1(m0_oper0_rdata_int[23]),.B0I2(NET_117),.B0I3(m1_oper1_rdata_int[23]),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[29]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_44),.T0I1(NET_117),.T0I2(m0_oper0_rdata_int[17]),.T0I3(m1_oper1_rdata_int[17]),.TB0S(GND),.B0Z(NET_455),.C0Z(NET_347),.Q0Z(tcdm_result_p0[29]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[23]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[23]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010101000000000),.B2I0(NET_346),.B2I1(tcdm_rdata_p0_int[17]),.B2I2(NET_124),.B2I3(NET_347),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[28]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_346),.T2I1(tcdm_rdata_p0_int[17]),.T2I2(NET_124),.T2I3(NET_347),.TB2S(NET_348),.C2Z(NET_330),.Q2Z(tcdm_result_p0[28]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010101000000000),.B3I0(NET_454),.B3I1(tcdm_rdata_p0_int[23]),.B3I2(NET_124),.B3I3(NET_455),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[19]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(NET_124),.T3I1(NET_455),.T3I2(NET_454),.T3I3(tcdm_rdata_p0_int[23]),.TB3S(NET_456),.C3Z(NET_439),.Q3Z(tcdm_result_p0[19]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_N12_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B0I0(tcdm_rdata_p1_int[22]),.B0I1(NET_110_CAND3_TLSBR_14_tpGCLKBUF),.B0I2(tcdm_rdata_p3_int[22]),.B0I3(NET_125_CAND4_TLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p1_int[22]),.T0I1(NET_110_CAND3_TLSBR_14_tpGCLKBUF),.T0I2(tcdm_rdata_p3_int[22]),.T0I3(NET_125_CAND4_TLSBR_14_tpGCLKBUF),.TB0S(NET_10),.C0Z(NET_435),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N12_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(tcdm_result_p1[22]),.B1I1(NET_89),.B1I2(NET_101),.B1I3(tcdm_result_p0[22]),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[18]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_101),.T1I1(tcdm_result_p0[22]),.T1I2(tcdm_result_p1[22]),.T1I3(NET_89),.TB1S(NET_15),.C1Z(NET_429),.Q1Z(tcdm_result_p1[18]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N12_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_101),.B2I1(tcdm_result_p0[18]),.B2I2(tcdm_result_p1[18]),.B2I3(NET_89),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[22]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_101),.T2I1(tcdm_result_p0[18]),.T2I2(tcdm_result_p1[18]),.T2I3(NET_89),.TB2S(NET_15),.C2Z(NET_357),.Q2Z(tcdm_result_p1[22]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N12_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B3I0(tcdm_result_p1[19]),.B3I1(NET_89),.B3I2(NET_101),.B3I3(tcdm_result_p0[19]),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[19]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(NET_101),.T3I1(tcdm_result_p0[19]),.T3I2(tcdm_result_p1[19]),.T3I3(NET_89),.TB3S(NET_15),.C3Z(NET_376),.Q3Z(tcdm_result_p1[19]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_N13_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_101),.B0I1(NET_89),.B0I2(tcdm_result_p0[23]),.B0I3(tcdm_result_p1[23]),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[22]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_101),.T0I1(NET_89),.T0I2(tcdm_result_p0[23]),.T0I3(tcdm_result_p1[23]),.TB0S(NET_15),.C0Z(NET_447),.Q0Z(tcdm_result_p3[22]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N13_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B1I0(tcdm_rdata_p1_int[23]),.B1I1(NET_110_CAND3_TLSBR_14_tpGCLKBUF),.B1I2(tcdm_rdata_p3_int[23]),.B1I3(NET_125_CAND4_TLSBR_14_tpGCLKBUF),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[23]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p3_int[23]),.T1I1(NET_125_CAND4_TLSBR_14_tpGCLKBUF),.T1I2(tcdm_rdata_p1_int[23]),.T1I3(NET_110_CAND3_TLSBR_14_tpGCLKBUF),.TB1S(NET_10),.C1Z(NET_453),.Q1Z(tcdm_result_p1[23]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N13_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B2I0(tcdm_result_p0[29]),.B2I1(NET_89),.B2I2(tcdm_result_p1[29]),.B2I3(NET_101),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[23]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p0[29]),.T2I1(NET_89),.T2I2(tcdm_result_p1[29]),.T2I3(NET_101),.TB2S(NET_15),.C2Z(NET_575),.Q2Z(tcdm_result_p3[23]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N13_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B3I0(tcdm_result_p1[28]),.B3I1(NET_101),.B3I2(tcdm_result_p0[28]),.B3I3(NET_89),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[18]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p0[28]),.T3I1(NET_89),.T3I2(tcdm_result_p1[28]),.T3I3(NET_101),.TB3S(NET_15),.C3Z(NET_557),.Q3Z(tcdm_result_p3[18]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_N14_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B0I0(tcdm_rdata_p1_int[28]),.B0I1(NET_125_CAND4_TLSBR_14_tpGCLKBUF),.B0I2(NET_110_CAND3_TLSBR_14_tpGCLKBUF),.B0I3(tcdm_rdata_p3_int[28]),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[28]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p1_int[28]),.T0I1(NET_125_CAND4_TLSBR_14_tpGCLKBUF),.T0I2(NET_110_CAND3_TLSBR_14_tpGCLKBUF),.T0I3(tcdm_rdata_p3_int[28]),.TB0S(NET_10),.C0Z(NET_563),.Q0Z(tcdm_result_p3[28]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N14_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(NET_125_CAND4_TLSBR_14_tpGCLKBUF),.B1I1(tcdm_rdata_p3_int[19]),.B1I2(tcdm_rdata_p1_int[19]),.B1I3(NET_110_CAND3_TLSBR_14_tpGCLKBUF),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[29]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p1_int[19]),.T1I1(NET_110_CAND3_TLSBR_14_tpGCLKBUF),.T1I2(NET_125_CAND4_TLSBR_14_tpGCLKBUF),.T1I3(tcdm_rdata_p3_int[19]),.TB1S(NET_10),.C1Z(NET_382),.Q1Z(tcdm_result_p3[29]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000010),.B2I0(lint_ADDR_int[7]),.B2I1(apb_fsm[0]),.B2I2(lint_ADDR_int[8]),.B2I3(lint_ADDR_int[11]),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[28]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[7]),.T2I1(apb_fsm[0]),.T2I2(lint_ADDR_int[8]),.T2I3(lint_ADDR_int[11]),.TB2S(lint_ADDR_int[2]),.C2Z(NET_101),.Q2Z(tcdm_result_p1[28]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N14_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B3I0(tcdm_rdata_p1_int[29]),.B3I1(tcdm_rdata_p3_int[29]),.B3I2(NET_110_CAND3_TLSBR_14_tpGCLKBUF),.B3I3(NET_125_CAND4_TLSBR_14_tpGCLKBUF),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[29]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(NET_110_CAND3_TLSBR_14_tpGCLKBUF),.T3I1(NET_125_CAND4_TLSBR_14_tpGCLKBUF),.T3I2(tcdm_rdata_p1_int[29]),.T3I3(tcdm_rdata_p3_int[29]),.TB3S(NET_10),.C3Z(NET_581),.Q3Z(tcdm_result_p1[29]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_N15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_75),.B0I1(NET_149),.B0I2(NET_71),.B0I3(NET_77),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_75),.T0I1(NET_149),.T0I2(NET_71),.T0I3(NET_77),.TB0S(NET_150),.C0Z(NET_147),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N15_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[0]),.T1I1(lint_ADDR_int[1]),.T1I2(GND),.T1I3(lint_ADDR_int[9]),.TB1S(GND),.C1Z(NET_71),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_N15_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000001000),.B2I0(NET_77),.B2I1(NET_69),.B2I2(GND),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[5]),.T2I1(GND),.T2I2(GND),.T2I3(lint_ADDR_int[7]),.TB2S(GND),.B2Z(NET_133),.C2Z(NET_75),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_N15_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[19]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[13]),.T3I1(GND),.T3I2(lint_ADDR_int[10]),.T3I3(lint_ADDR_int[4]),.TB3S(GND),.C3Z(NET_150),.Q3Z(tcdm_result_p3[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_N16_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000001000000000),.B0I0(NET_69),.B0I1(lint_ADDR_int[4]),.B0I2(lint_ADDR_int[5]),.B0I3(NET_77),.T0I0(lint_ADDR_int[11]),.T0I1(GND),.T0I2(GND),.T0I3(lint_ADDR_int[6]),.TB0S(GND),.B0Z(NET_173),.C0Z(NET_77),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_N16_1 (.tFragBitInfo(16'b0000000001011101),.bFragBitInfo(16'b0001001100010011),.B1I0(NET_75),.B1I1(NET_622),.B1I2(NET_77),.B1I3(lint_ADDR_int[4]),.T1I0(NET_77),.T1I1(lint_ADDR_int[4]),.T1I2(NET_75),.T1I3(NET_622),.TB1S(lint_ADDR_int[5]),.C1Z(NET_754),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_N16_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0010000000000000),.B2I0(NET_69),.B2I1(GND),.B2I2(NET_75),.B2I3(NET_77),.T2I0(NET_69),.T2I1(NET_131),.T2I2(NET_622),.T2I3(NET_65),.TB2S(GND),.B2Z(NET_66),.C2Z(nx60509z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_N16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000100),.B3I0(lint_ADDR_int[7]),.B3I1(lint_ADDR_int[6]),.B3I2(lint_ADDR_int[11]),.B3I3(lint_ADDR_int[4]),.T3I0(lint_ADDR_int[11]),.T3I1(lint_ADDR_int[4]),.T3I2(lint_ADDR_int[7]),.T3I3(lint_ADDR_int[6]),.TB3S(lint_ADDR_int[5]),.C3Z(NET_622),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_N17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N17_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_172),.T1I1(GND),.T1I2(NET_66),.T1I3(GND),.TB1S(GND),.C1Z(nx23147z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_N17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_65),.B2I1(NET_131),.B2I2(GND),.B2I3(lint_ADDR_int[4]),.B2Z(NET_172),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N18_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.B1I0(m1_ram_control[25]),.B1I1(NET_17_CAND2_BLSTR_14_tpGCLKBUF),.B1I2(m1_m1_control[25]),.B1I3(NET_28_CAND5_BLSTR_14_tpGCLKBUF),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx49871z1_CAND3_BLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_control[25]),.T1I1(NET_28_CAND5_BLSTR_14_tpGCLKBUF),.T1I2(m1_ram_control[25]),.T1I3(NET_17_CAND2_BLSTR_14_tpGCLKBUF),.TB1S(NET_505),.C1Z(NET_503),.Q1Z(m1_ram_control[25]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m1_m1_control[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_sat_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N19_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.B1I0(m1_ram_control[16]),.B1I1(NET_28_CAND5_BLSTR_14_tpGCLKBUF),.B1I2(m1_m1_rnd_dup_0),.B1I3(NET_17_CAND2_BLSTR_14_tpGCLKBUF),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx49871z1_CAND3_BLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_rnd_dup_0),.T1I1(NET_17_CAND2_BLSTR_14_tpGCLKBUF),.T1I2(m1_ram_control[16]),.T1I3(NET_28_CAND5_BLSTR_14_tpGCLKBUF),.TB1S(NET_321),.C1Z(NET_319),.Q1Z(m1_ram_control[16]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N19_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.B2I0(m1_m1_reset_dup_0),.B2I1(NET_17_CAND2_BLSTR_14_tpGCLKBUF),.B2I2(m1_ram_control[31]),.B2I3(NET_28_CAND5_BLSTR_14_tpGCLKBUF),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx49871z1_CAND3_BLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T2I0(m1_m1_reset_dup_0),.T2I1(NET_17_CAND2_BLSTR_14_tpGCLKBUF),.T2I2(m1_ram_control[31]),.T2I3(NET_28_CAND5_BLSTR_14_tpGCLKBUF),.TB2S(NET_612),.C2Z(NET_610),.Q2Z(m1_ram_control[31]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_reset_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m1_m1_rnd_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m1_m1_osel_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[6]),.Q0EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_waddr_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[8]),.Q1EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[9]),.Q2EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_waddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[8]),.Q3EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_waddr_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(NET_762),.Q0EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_we_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[11]),.Q1EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[2]),.Q2EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_waddr_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[3]),.Q3EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_waddr_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N32_0 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0000000000101010),.B0I0(NET_748),.B0I1(m1_coef_rdata_int[27]),.B0I2(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.B0I3(m1_oper1_rdata_int[27]),.CD0S(VCC),.Q0DI(lint_ADDR_int[9]),.Q0EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_748),.T0I1(m1_coef_rdata_int[27]),.T0I2(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.T0I3(m1_oper1_rdata_int[27]),.TB0S(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.C0Z(NET_749),.Q0Z(m1_coef_raddr_dup_0[9]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N32_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[7]),.Q1EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.T1I1(m1_oper1_rdata_int[1]),.T1I2(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.T1I3(m1_coef_rdata_int[1]),.TB1S(GND),.C1Z(NET_39),.Q1Z(m1_coef_waddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N32_2 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0000000000101010),.B2I0(NET_742),.B2I1(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.B2I2(m1_coef_rdata_int[16]),.B2I3(m1_oper1_rdata_int[16]),.CD2S(VCC),.Q2DI(lint_ADDR_int[1]),.Q2EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_742),.T2I1(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.T2I2(m1_coef_rdata_int[16]),.T2I3(m1_oper1_rdata_int[16]),.TB2S(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.C2Z(NET_743),.Q2Z(m1_coef_waddr_dup_0[1]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N32_3 (.tFragBitInfo(16'b0011111100000000),.bFragBitInfo(16'b0000010000001100),.B3I0(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.B3I1(NET_746),.B3I2(m1_oper1_rdata_int[25]),.B3I3(m1_coef_rdata_int[25]),.CD3S(VCC),.Q3DI(lint_ADDR_int[5]),.Q3EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(m1_oper1_rdata_int[25]),.T3I1(m1_coef_rdata_int[25]),.T3I2(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.T3I3(NET_746),.TB3S(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.C3Z(NET_747),.Q3Z(m1_coef_waddr_dup_0[5]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_O1_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[4]),.Q0EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.T0I0(m0_coef_rdata_int[31]),.T0I1(NET_41_CAND4_TLSTR_15_tpGCLKBUF),.T0I2(NET_46_CAND3_TLSTR_15_tpGCLKBUF),.T0I3(m0_oper1_rdata_int[31]),.TB0S(GND),.C0Z(NET_615),.Q0Z(m0_coef_raddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O1_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[1]),.Q1EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.T1I0(NET_46_CAND3_TLSTR_15_tpGCLKBUF),.T1I1(NET_41_CAND4_TLSTR_15_tpGCLKBUF),.T1I2(m0_coef_rdata_int[20]),.T1I3(m0_oper1_rdata_int[20]),.TB1S(GND),.C1Z(NET_398),.Q1Z(m0_coef_raddr_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_O1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[0]),.Q2EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_raddr_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O1_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.T3I0(m0_coef_rdata_int[19]),.T3I1(m0_oper1_rdata_int[19]),.T3I2(NET_46_CAND3_TLSTR_15_tpGCLKBUF),.T3I3(NET_41_CAND4_TLSTR_15_tpGCLKBUF),.C3Z(NET_385),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[2]),.Q0EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_raddr_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[5]),.Q1EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_raddr_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[3]),.Q2EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_raddr_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[6]),.Q3EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_raddr_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[7]),.Q1EN(nx32231z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_raddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O7_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p0_int[4]),.T0I1(NET_62),.T0I2(m0_m1_outsel_dup_0[4]),.T0I3(NET_63),.TB0S(GND),.C0Z(NET_682),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_outsel_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O9_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000100),.B0I0(lint_ADDR_int[3]),.B0I1(lint_ADDR_int[4]),.B0I2(lint_ADDR_int[2]),.B0I3(GND),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(NET_65),.T0I1(NET_133),.T0I2(NET_531),.T0I3(NET_139),.TB0S(GND),.B0Z(NET_138),.Q0Z(m0_m1_clken_dup_0),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O9_1 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[3]),.T1I1(lint_ADDR_int[4]),.T1I2(lint_ADDR_int[2]),.T1I3(GND),.TB1S(GND),.C1Z(NET_531),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_O9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O9_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_65),.T3I1(NET_133),.T3I2(NET_138),.T3I3(NET_139),.TB3S(GND),.Q3Z(m0_m0_clken_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_O10_0 (.tFragBitInfo(16'b1010000000000000),.bFragBitInfo(16'b0010000000000000),.B0I0(NET_753),.B0I1(m0_oper0_rdata_int[31]),.B0I2(NET_615),.B0I3(NET_614),.T0I0(NET_753),.T0I1(m0_oper0_rdata_int[31]),.T0I2(NET_615),.T0I3(NET_614),.TB0S(NET_117),.C0Z(NET_606),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_O10_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[5]),.T1I1(lint_ADDR_int[3]),.T1I2(lint_ADDR_int[6]),.T1I3(lint_ADDR_int[4]),.C1Z(NET_15),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O10_2 (.tFragBitInfo(16'b1000100000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_597),.B2I1(NET_751),.B2I2(m0_oper0_rdata_int[30]),.B2I3(NET_596),.T2I0(NET_597),.T2I1(NET_751),.T2I2(m0_oper0_rdata_int[30]),.T2I3(NET_596),.TB2S(NET_117),.C2Z(NET_588),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_O10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000011000000),.B1I0(NET_124),.B1I1(NET_528),.B1I2(NET_529),.B1I3(tcdm_rdata_p0_int[26]),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[24]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(NET_529),.T1I1(tcdm_rdata_p0_int[26]),.T1I2(NET_124),.T1I3(NET_528),.TB1S(NET_530),.C1Z(NET_513),.Q1Z(tcdm_result_p0[24]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_O11_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_117),.B2I1(NET_44),.B2I2(m0_oper0_rdata_int[26]),.B2I3(m1_oper1_rdata_int[26]),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_rdata_int[24]),.T2I1(NET_44),.T2I2(NET_117),.T2I3(m0_oper0_rdata_int[24]),.TB2S(GND),.B2Z(NET_529),.C2Z(NET_494),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_O11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100110000000000),.B3I0(NET_124),.B3I1(NET_493),.B3I2(tcdm_rdata_p0_int[24]),.B3I3(NET_494),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[21]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p0_int[24]),.T3I1(NET_494),.T3I2(NET_124),.T3I3(NET_493),.TB3S(NET_495),.C3Z(NET_478),.Q3Z(tcdm_result_p0[21]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_O12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[17]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p1[17]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O12_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B1I0(NET_110_CAND3_TLSBR_15_tpGCLKBUF),.B1I1(NET_125_CAND4_TLSBR_15_tpGCLKBUF),.B1I2(tcdm_rdata_p1_int[17]),.B1I3(tcdm_rdata_p3_int[17]),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[17]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p1_int[17]),.T1I1(tcdm_rdata_p3_int[17]),.T1I2(NET_110_CAND3_TLSBR_15_tpGCLKBUF),.T1I3(NET_125_CAND4_TLSBR_15_tpGCLKBUF),.TB1S(NET_10),.C1Z(NET_345),.Q1Z(tcdm_result_p0[17]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_O12_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B2I0(tcdm_result_p0[21]),.B2I1(NET_101),.B2I2(NET_89),.B2I3(tcdm_result_p1[21]),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p0[21]),.T2I1(NET_101),.T2I2(NET_89),.T2I3(tcdm_result_p1[21]),.TB2S(NET_15),.C2Z(NET_411),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_O12_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B3I0(tcdm_result_p0[17]),.B3I1(NET_89),.B3I2(tcdm_result_p1[17]),.B3I3(NET_101),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[21]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p1[17]),.T3I1(NET_101),.T3I2(tcdm_result_p0[17]),.T3I3(NET_89),.TB3S(NET_15),.C3Z(NET_339),.Q3Z(tcdm_result_p1[21]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_O13_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_101),.B0I1(NET_89),.B0I2(tcdm_result_p0[24]),.B0I3(tcdm_result_p1[24]),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[26]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(NET_101),.T0I1(NET_89),.T0I2(tcdm_result_p0[24]),.T0I3(tcdm_result_p1[24]),.TB0S(NET_15),.C0Z(NET_486),.Q0Z(tcdm_result_p1[26]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O13_1 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[26]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(NET_89),.T1I2(NET_7),.T1I3(GND),.C1Z(NET_82),.Q1Z(tcdm_result_p0[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O13_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_101),.B2I1(NET_89),.B2I2(tcdm_result_p0[26]),.B2I3(tcdm_result_p1[26]),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[17]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_101),.T2I1(NET_89),.T2I2(tcdm_result_p0[26]),.T2I3(tcdm_result_p1[26]),.TB2S(NET_15),.C2Z(NET_521),.Q2Z(tcdm_result_p3[17]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O13_3 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_101),.T3I1(GND),.T3I2(NET_7),.T3I3(GND),.C3Z(NET_99),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O14_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(tcdm_result_p3[7]),.B0I1(tcdm_result_p1[7]),.B0I2(NET_99),.B0I3(NET_100),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[7]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p1[2]),.T0I1(NET_99),.T0I2(tcdm_result_p3[2]),.T0I3(NET_100),.TB0S(GND),.B0Z(NET_463),.C0Z(NET_711),.Q0Z(tcdm_result_p1[7]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O14_1 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[2]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(NET_15),.T1I2(GND),.T1I3(NET_101),.C1Z(NET_100),.Q1Z(tcdm_result_p1[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O14_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_125_CAND4_TLSBR_15_tpGCLKBUF),.B2I1(NET_110_CAND3_TLSBR_15_tpGCLKBUF),.B2I2(tcdm_rdata_p3_int[2]),.B2I3(tcdm_rdata_p1_int[2]),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[26]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_125_CAND4_TLSBR_15_tpGCLKBUF),.T2I1(NET_110_CAND3_TLSBR_15_tpGCLKBUF),.T2I2(tcdm_rdata_p3_int[2]),.T2I3(tcdm_rdata_p1_int[2]),.TB2S(NET_10),.C2Z(NET_725),.Q2Z(tcdm_result_p3[26]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O14_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B3I0(tcdm_rdata_p1_int[26]),.B3I1(tcdm_rdata_p3_int[26]),.B3I2(NET_125_CAND4_TLSBR_15_tpGCLKBUF),.B3I3(NET_110_CAND3_TLSBR_15_tpGCLKBUF),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[2]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_125_CAND4_TLSBR_15_tpGCLKBUF),.T3I1(NET_110_CAND3_TLSBR_15_tpGCLKBUF),.T3I2(tcdm_rdata_p1_int[26]),.T3I3(tcdm_rdata_p3_int[26]),.TB3S(NET_10),.C3Z(NET_527),.Q3Z(tcdm_result_p3[2]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_O15_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_99),.B0I1(tcdm_result_p3[12]),.B0I2(tcdm_result_p1[12]),.B0I3(NET_100),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[6]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(NET_99),.T0I1(tcdm_result_p1[0]),.T0I2(tcdm_result_p3[0]),.T0I3(NET_100),.TB0S(GND),.B0Z(NET_219),.C0Z(NET_91),.Q0Z(tcdm_result_p3[6]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O15_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B1I0(tcdm_rdata_p1_int[6]),.B1I1(NET_125_CAND4_TLSBR_15_tpGCLKBUF),.B1I2(NET_110_CAND3_TLSBR_15_tpGCLKBUF),.B1I3(tcdm_rdata_p3_int[6]),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[6]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(NET_110_CAND3_TLSBR_15_tpGCLKBUF),.T1I1(tcdm_rdata_p3_int[6]),.T1I2(tcdm_rdata_p1_int[6]),.T1I3(NET_125_CAND4_TLSBR_15_tpGCLKBUF),.TB1S(NET_10),.C1Z(NET_643),.Q1Z(tcdm_result_p1[6]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_O15_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_125_CAND4_TLSBR_15_tpGCLKBUF),.B2I1(tcdm_rdata_p3_int[0]),.B2I2(tcdm_rdata_p1_int[0]),.B2I3(NET_110_CAND3_TLSBR_15_tpGCLKBUF),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[0]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_125_CAND4_TLSBR_15_tpGCLKBUF),.T2I1(tcdm_rdata_p3_int[0]),.T2I2(tcdm_rdata_p1_int[0]),.T2I3(NET_110_CAND3_TLSBR_15_tpGCLKBUF),.TB2S(NET_10),.C2Z(NET_130),.Q2Z(tcdm_result_p1[0]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O15_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[0]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_99),.T3I1(tcdm_result_p3[6]),.T3I2(tcdm_result_p1[6]),.T3I3(NET_100),.C3Z(NET_629),.Q3Z(tcdm_result_p3[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000010000),.B0I0(GND),.B0I1(GND),.B0I2(lint_ADDR_int[5]),.B0I3(lint_ADDR_int[7]),.B0Z(NET_139),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O16_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_10),.T1I1(tcdm_rdata_p1_int[31]),.T1I2(NET_15),.T1I3(GND),.TB1S(GND),.C1Z(NET_612),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_O16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000010),.B2I0(lint_ADDR_int[8]),.B2I1(GND),.B2I2(GND),.B2I3(apb_fsm[0]),.B2Z(NET_19),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O16_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_10),.T3I1(GND),.T3I2(NET_15),.T3I3(tcdm_rdata_p1_int[16]),.TB3S(GND),.C3Z(NET_321),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_O17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001000),.B0I0(lint_ADDR_int[3]),.B0I1(lint_ADDR_int[4]),.B0I2(lint_ADDR_int[2]),.B0I3(GND),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.B0Z(NET_646),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O17_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_139),.T2I1(NET_133),.T2I2(GND),.T2I3(NET_172),.TB2S(GND),.Q2Z(m1_m1_clken_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_O17_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_139),.T3I1(NET_133),.T3I2(NET_646),.T3I3(NET_65),.TB3S(GND),.Q3Z(m1_m0_clken_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_O31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[3]),.Q0EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_raddr_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[6]),.Q1EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_oper1_rdata_int[4]),.B2I1(NET_44_CAND4_BLSBR_15_tpGCLKBUF),.B2I2(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.B2I3(m1_coef_rdata_int[4]),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.B2Z(NET_677),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[2]),.Q3EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_raddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O32_0 (.tFragBitInfo(16'b0000110011001100),.bFragBitInfo(16'b0000010001000100),.B0I0(m1_oper1_rdata_int[30]),.B0I1(NET_750),.B0I2(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.B0I3(m1_coef_rdata_int[30]),.CD0S(VCC),.Q0DI(lint_ADDR_int[1]),.Q0EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_rdata_int[30]),.T0I1(NET_750),.T0I2(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.T0I3(m1_coef_rdata_int[30]),.TB0S(NET_44_CAND4_BLSBR_15_tpGCLKBUF),.C0Z(NET_751),.Q0Z(m1_coef_raddr_dup_0[1]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O32_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(NET_44_CAND4_BLSBR_15_tpGCLKBUF),.T1I1(m1_oper1_rdata_int[8]),.T1I2(m1_coef_rdata_int[8]),.T1I3(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.C1Z(NET_283),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O32_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[4]),.Q2EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_44_CAND4_BLSBR_15_tpGCLKBUF),.T2I1(m1_coef_rdata_int[5]),.T2I2(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.T2I3(m1_oper1_rdata_int[5]),.TB2S(GND),.C2Z(NET_657),.Q2Z(m1_coef_raddr_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O32_3 (.tFragBitInfo(16'b0100010011001100),.bFragBitInfo(16'b0001010100000000),.B3I0(m1_oper1_rdata_int[31]),.B3I1(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.B3I2(m1_coef_rdata_int[31]),.B3I3(NET_752),.CD3S(VCC),.Q3DI(lint_ADDR_int[7]),.Q3EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(m1_coef_rdata_int[31]),.T3I1(NET_752),.T3I2(m1_oper1_rdata_int[31]),.T3I3(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.TB3S(NET_44_CAND4_BLSBR_15_tpGCLKBUF),.C3Z(NET_753),.Q3Z(m1_coef_raddr_dup_0[7]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_P1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_41_CAND4_TLSTR_16_tpGCLKBUF),.B0I1(m0_coef_rdata_int[18]),.B0I2(NET_46_CAND3_TLSTR_16_tpGCLKBUF),.B0I3(m0_oper1_rdata_int[18]),.B0Z(NET_366),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P1_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_oper1_rdata_int[30]),.T1I1(NET_41_CAND4_TLSTR_16_tpGCLKBUF),.T1I2(m0_coef_rdata_int[30]),.T1I3(NET_46_CAND3_TLSTR_16_tpGCLKBUF),.C1Z(NET_597),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_P1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_41_CAND4_TLSTR_16_tpGCLKBUF),.B2I1(m0_coef_rdata_int[17]),.B2I2(NET_46_CAND3_TLSTR_16_tpGCLKBUF),.B2I3(m0_oper1_rdata_int[17]),.B2Z(NET_348),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P1_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_41_CAND4_TLSTR_16_tpGCLKBUF),.T3I1(NET_46_CAND3_TLSTR_16_tpGCLKBUF),.T3I2(m0_oper1_rdata_int[24]),.T3I3(m0_coef_rdata_int[24]),.C3Z(NET_495),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_outsel_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P7_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p0_int[1]),.T1I1(NET_63),.T1I2(NET_62),.T1I3(m0_m1_outsel_dup_0[1]),.TB1S(GND),.C1Z(NET_54),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_P7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_mode_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_csel_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m0_m1_csel_dup_0),.B2I1(NET_63),.B2I2(NET_62),.B2I3(tcdm_rdata_p0_int[15]),.B2Z(NET_307),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P10_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_51),.B0I1(NET_63),.B0I2(tcdm_result_p3[25]),.B0I3(m0_m1_control[25]),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(NET_51),.T0I1(NET_63),.T0I2(tcdm_result_p3[27]),.T0I3(m0_m1_control[27]),.TB0S(GND),.B0Z(NET_507),.C0Z(NET_543),.Q0Z(m0_m1_control[27]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[20]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_control[20]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P10_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T3I0(NET_51),.T3I1(tcdm_result_p3[20]),.T3I2(m0_m1_control[20]),.T3I3(NET_63),.C3Z(NET_397),.Q3Z(m0_m1_control[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P12_0 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[27]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[6]),.T0I1(lint_ADDR_int[5]),.T0I2(NET_146),.T0I3(NET_145),.TB0S(GND),.C0Z(nx49871z1),.Q0Z(tcdm_result_p3[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[20]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[20]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P13_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B0I0(tcdm_rdata_p1_int[24]),.B0I1(tcdm_rdata_p3_int[24]),.B0I2(NET_110_CAND3_TLSBR_16_tpGCLKBUF),.B0I3(NET_125_CAND4_TLSBR_16_tpGCLKBUF),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[24]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p1_int[24]),.T0I1(tcdm_rdata_p3_int[24]),.T0I2(NET_110_CAND3_TLSBR_16_tpGCLKBUF),.T0I3(NET_125_CAND4_TLSBR_16_tpGCLKBUF),.TB0S(NET_10),.C0Z(NET_492),.Q0Z(tcdm_result_p1[24]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[25]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p3[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B2I0(lint_ADDR_int[6]),.B2I1(lint_ADDR_int[4]),.B2I2(lint_ADDR_int[5]),.B2I3(lint_ADDR_int[11]),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[24]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[6]),.T2I1(lint_ADDR_int[4]),.T2I2(lint_ADDR_int[5]),.T2I3(lint_ADDR_int[11]),.TB2S(lint_ADDR_int[3]),.C2Z(NET_110),.Q2Z(tcdm_result_p3[24]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_P13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P14_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(tcdm_rdata_p1_int[7]),.B0I1(NET_110_CAND3_TLSBR_16_tpGCLKBUF),.B0I2(NET_125_CAND4_TLSBR_16_tpGCLKBUF),.B0I3(tcdm_rdata_p3_int[7]),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[21]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p1_int[7]),.T0I1(NET_110_CAND3_TLSBR_16_tpGCLKBUF),.T0I2(NET_125_CAND4_TLSBR_16_tpGCLKBUF),.T0I3(tcdm_rdata_p3_int[7]),.TB0S(NET_10),.C0Z(NET_477),.Q0Z(tcdm_result_p3[21]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P14_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[7]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T1I0(NET_10),.T1I1(NET_15),.T1I2(GND),.T1I3(tcdm_rdata_p1_int[20]),.TB1S(GND),.C1Z(NET_395),.Q1Z(tcdm_result_p3[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_P14_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_110_CAND3_TLSBR_16_tpGCLKBUF),.B2I1(tcdm_rdata_p1_int[21]),.B2I2(NET_125_CAND4_TLSBR_16_tpGCLKBUF),.B2I3(tcdm_rdata_p3_int[21]),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T2I0(NET_110_CAND3_TLSBR_16_tpGCLKBUF),.T2I1(tcdm_rdata_p1_int[21]),.T2I2(NET_125_CAND4_TLSBR_16_tpGCLKBUF),.T2I3(tcdm_rdata_p3_int[21]),.TB2S(NET_10),.C2Z(NET_417),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_P14_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p1_int[30]),.T3I1(NET_15),.T3I2(NET_10),.T3I3(GND),.TB3S(GND),.C3Z(NET_594),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_P15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P15_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(tcdm_rdata_p1_int[12]),.B1I1(tcdm_rdata_p3_int[12]),.B1I2(NET_125_CAND4_TLSBR_16_tpGCLKBUF),.B1I3(NET_110_CAND3_TLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T1I0(NET_125_CAND4_TLSBR_16_tpGCLKBUF),.T1I1(NET_110_CAND3_TLSBR_16_tpGCLKBUF),.T1I2(tcdm_rdata_p1_int[12]),.T1I3(tcdm_rdata_p3_int[12]),.TB1S(NET_10),.C1Z(NET_233),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_P15_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.B2I0(lint_ADDR_int[3]),.B2I1(lint_ADDR_int[4]),.B2I2(lint_ADDR_int[5]),.B2I3(lint_ADDR_int[11]),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[12]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[3]),.T2I1(lint_ADDR_int[4]),.T2I2(lint_ADDR_int[5]),.T2I3(lint_ADDR_int[11]),.TB2S(lint_ADDR_int[6]),.C2Z(NET_125),.Q2Z(tcdm_result_p3[12]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_P15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[12]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p1[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000010000000000),.B0I0(GND),.B0I1(NET_14),.B0I2(GND),.B0I3(NET_15),.B0Z(NET_13),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P16_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(tcdm_rdata_p1_int[25]),.T1I1(NET_10),.T1I2(GND),.T1I3(NET_15),.TB1S(GND),.C1Z(NET_505),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_P16_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(tcdm_rdata_p1_int[27]),.T2I1(NET_10),.T2I2(GND),.T2I3(NET_15),.TB2S(GND),.C2Z(NET_541),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_P16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[10]),.Q1EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[5]),.Q2EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_raddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[0]),.Q3EN(nx14650z1),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_raddr_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m0_oper1_rdata_int[26]),.B0I1(NET_46),.B0I2(NET_41),.B0I3(m0_coef_rdata_int[26]),.B0Z(NET_530),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q1_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_oper1_rdata_int[25]),.T1I1(NET_46),.T1I2(m0_coef_rdata_int[25]),.T1I3(NET_41),.C1Z(NET_508),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Q1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(m0_coef_rdata_int[27]),.B2I1(NET_46),.B2I2(m0_oper1_rdata_int[27]),.B2I3(NET_41),.B2Z(NET_544),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q1_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m0_oper1_rdata_int[21]),.T3I1(m0_coef_rdata_int[21]),.T3I2(NET_46),.T3I3(NET_41),.C3Z(NET_420),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_Q2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q2_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_46),.T1I1(NET_41),.T1I2(m0_oper1_rdata_int[23]),.T1I3(m0_coef_rdata_int[23]),.C1Z(NET_456),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Q2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.Q2Z(m0_m1_reset_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.Q3Z(m0_m1_outsel_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.Q1Z(m0_m1_outsel_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q7_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.T2I0(tcdm_rdata_p0_int[3]),.T2I1(NET_62),.T2I2(m0_m1_outsel_dup_0[3]),.T2I3(NET_63),.TB2S(GND),.C2Z(NET_701),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_Q7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.Q1Z(m0_m1_sat_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.Q2Z(m0_m1_tc_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0),.QST(GND),.Q3Z(m0_m1_rnd_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q10_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T0I0(NET_63),.T0I1(tcdm_result_p3[30]),.T0I2(m0_m1_control[30]),.T0I3(NET_51),.TB0S(GND),.C0Z(NET_596),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q10_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_63),.B2I1(NET_51),.B2I2(m0_m1_rnd_dup_0),.B2I3(tcdm_result_p3[16]),.CD2S(VCC),.Q2DI(lint_WDATA_int[30]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T2I0(NET_63),.T2I1(NET_51),.T2I2(m0_m1_reset_dup_0),.T2I3(tcdm_result_p3[31]),.TB2S(GND),.B2Z(NET_324),.C2Z(NET_614),.Q2Z(m0_m1_control[30]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_Q10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[3]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[31]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p3[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[30]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[30]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[16]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p3[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q13_0 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[16]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[11]),.T0I1(GND),.T0I2(apb_fsm[0]),.T0I3(lint_ADDR_int[8]),.TB0S(GND),.C0Z(NET_87),.Q0Z(tcdm_result_p0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q13_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[27]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T1I0(NET_50_CAND4_TRSBL_17_tpGCLKBUF),.T1I1(NET_62),.T1I2(tcdm_result_p1[16]),.T1I3(tcdm_rdata_p0_int[16]),.TB1S(GND),.C1Z(NET_316),.Q1Z(tcdm_result_p0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_Q13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001000),.B2I0(NET_49),.B2I1(NET_7),.B2I2(GND),.B2I3(GND),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[27]),.Q2EN(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B2Z(NET_51),.Q2Z(tcdm_result_p1[27]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q13_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[16]),.Q3EN(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p1[27]),.T3I1(NET_62),.T3I2(tcdm_rdata_p0_int[27]),.T3I3(NET_50_CAND4_TRSBL_17_tpGCLKBUF),.TB3S(GND),.C3Z(NET_536),.Q3Z(tcdm_result_p1[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Q14_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B0I0(tcdm_rdata_p0_int[20]),.B0I1(NET_62),.B0I2(tcdm_result_p1[20]),.B0I3(NET_50_CAND4_TRSBL_17_tpGCLKBUF),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[30]),.Q0EN(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p0_int[31]),.T0I1(NET_62),.T0I2(tcdm_result_p1[31]),.T0I3(NET_50_CAND4_TRSBL_17_tpGCLKBUF),.TB0S(GND),.B0Z(NET_390),.C0Z(NET_607),.Q0Z(tcdm_result_p1[30]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q14_1 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[20]),.Q1EN(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(NET_15),.T1I2(NET_49),.T1I3(GND),.C1Z(NET_50),.Q1Z(tcdm_result_p1[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Q14_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[31]),.Q2EN(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p1[30]),.T2I1(NET_62),.T2I2(tcdm_rdata_p0_int[30]),.T2I3(NET_50_CAND4_TRSBL_17_tpGCLKBUF),.TB2S(GND),.C2Z(NET_589),.Q2Z(tcdm_result_p1[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_Q14_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[25]),.Q3EN(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p0_int[25]),.T3I1(NET_62),.T3I2(tcdm_result_p1[25]),.T3I3(NET_50_CAND4_TRSBL_17_tpGCLKBUF),.TB3S(GND),.C3Z(NET_500),.Q3Z(tcdm_result_p1[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Q15_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_13),.B0I1(tcdm_rdata_p3_int[27]),.B0I2(NET_34),.B0I3(tcdm_result_p0[27]),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[20]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T0I0(NET_13),.T0I1(tcdm_result_p0[30]),.T0I2(NET_34),.T0I3(tcdm_rdata_p3_int[30]),.TB0S(GND),.B0Z(NET_547),.C0Z(NET_600),.Q0Z(tcdm_result_p0[20]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q15_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[25]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T1I0(NET_13),.T1I1(tcdm_result_p0[20]),.T1I2(NET_34),.T1I3(tcdm_rdata_p3_int[20]),.TB1S(GND),.C1Z(NET_401),.Q1Z(tcdm_result_p0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_Q15_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_13),.B2I1(tcdm_rdata_p3_int[25]),.B2I2(NET_34),.B2I3(tcdm_result_p0[25]),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[30]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T2I0(NET_13),.T2I1(tcdm_rdata_p3_int[16]),.T2I2(NET_34),.T2I3(tcdm_result_p0[16]),.TB2S(GND),.B2Z(NET_511),.C2Z(NET_328),.Q2Z(tcdm_result_p0[30]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_Q15_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[31]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T3I0(NET_13),.T3I1(tcdm_rdata_p3_int[31]),.T3I2(NET_34),.T3I3(tcdm_result_p0[31]),.TB3S(GND),.C3Z(NET_618),.Q3Z(tcdm_result_p0[31]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Q17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000010),.B0I0(lint_ADDR_int[7]),.B0I1(lint_ADDR_int[2]),.B0I2(apb_fsm[0]),.B0I3(lint_ADDR_int[8]),.B0Z(NET_14),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q17_1 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[7]),.T1I1(lint_ADDR_int[2]),.T1I2(apb_fsm[0]),.T1I3(lint_ADDR_int[8]),.C1Z(NET_49),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Q17_2 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'b0000000000000000),.T2I0(GND),.T2I1(lint_ADDR_int[2]),.T2I2(GND),.T2I3(NET_65),.TB2S(GND),.C2Z(NET_134),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_Q17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q18_0 (.tFragBitInfo(16'b0000000000000100),.bFragBitInfo(16'b0000000000000000),.T0I0(lint_ADDR_int[8]),.T0I1(lint_ADDR_int[2]),.T0I2(lint_ADDR_int[7]),.T0I3(apb_fsm[0]),.TB0S(GND),.C0Z(NET_10),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_Q18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R10_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_85),.B0I1(NET_86),.B0I2(m0_m1_dataout_int[0]),.B0I3(m1_ram_control[0]),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(NET_85),.T0I1(NET_86),.T0I2(m1_ram_control[12]),.T0I3(m0_m1_dataout_int[12]),.TB0S(GND),.B0Z(NET_84),.C0Z(NET_217),.Q0Z(m1_ram_control[0]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R10_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(NET_85),.T1I1(m0_m1_dataout_int[2]),.T1I2(m1_ram_control[2]),.T1I3(NET_86),.TB1S(GND),.C1Z(NET_709),.Q1Z(m1_ram_control[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_R10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.Q2Z(m1_ram_control[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R11_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(m0_m1_dataout_int[29]),.T0I1(m1_m1_dataout_int[29]),.T0I2(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.T0I3(NET_86),.TB0S(GND),.C0Z(NET_571),.Q0Z(m1_ram_control[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R11_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(NET_85),.T1I1(m1_ram_control[7]),.T1I2(m0_m1_dataout_int[7]),.T1I3(NET_86),.TB1S(GND),.C1Z(NET_461),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_R11_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(NET_86),.T2I1(m0_m1_dataout_int[26]),.T2I2(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.T2I3(m1_m1_dataout_int[26]),.TB2S(GND),.C2Z(NET_517),.Q2Z(m1_ram_control[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_R11_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T3I0(NET_85),.T3I1(m0_m1_dataout_int[6]),.T3I2(NET_86),.T3I3(m1_ram_control[6]),.C3Z(NET_627),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_R12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_82),.B0I1(m1_m1_dataout_int[7]),.B0I2(tcdm_result_p2[7]),.B0I3(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(NET_82),.T0I1(m1_m1_dataout_int[7]),.T0I2(tcdm_result_p2[7]),.T0I3(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.TB0S(NET_461),.C0Z(NET_459),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R12_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_dataout_int[28]),.T1I1(NET_86),.T1I2(m0_m1_dataout_int[28]),.T1I3(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.C1Z(NET_553),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_R12_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(NET_15),.T2I1(NET_87),.T2I2(lint_ADDR_int[2]),.T2I3(lint_ADDR_int[7]),.TB2S(GND),.C2Z(NET_86),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_R12_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[7]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T3I0(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.T3I1(m0_m1_dataout_int[24]),.T3I2(NET_86),.T3I3(m1_m1_dataout_int[24]),.TB3S(GND),.C3Z(NET_482),.Q3Z(tcdm_result_p2[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_R13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m1_m1_dataout_int[12]),.B0I1(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.B0I2(NET_82),.B0I3(tcdm_result_p2[12]),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[2]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(m1_m1_dataout_int[12]),.T0I1(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.T0I2(NET_82),.T0I3(tcdm_result_p2[12]),.TB0S(NET_217),.C0Z(NET_215),.Q0Z(tcdm_result_p2[2]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B1I0(NET_82),.B1I1(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.B1I2(m1_m1_dataout_int[2]),.B1I3(tcdm_result_p2[2]),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[0]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_dataout_int[2]),.T1I1(tcdm_result_p2[2]),.T1I2(NET_82),.T1I3(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.TB1S(NET_709),.C1Z(NET_707),.Q1Z(tcdm_result_p2[0]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_R13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.B2I1(m1_m1_dataout_int[0]),.B2I2(NET_82),.B2I3(tcdm_result_p2[0]),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[6]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.T2I1(m1_m1_dataout_int[0]),.T2I2(NET_82),.T2I3(tcdm_result_p2[0]),.TB2S(NET_84),.C2Z(NET_80),.Q2Z(tcdm_result_p2[6]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_R13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(NET_82),.B3I1(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.B3I2(tcdm_result_p2[6]),.B3I3(m1_m1_dataout_int[6]),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[12]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p2[6]),.T3I1(m1_m1_dataout_int[6]),.T3I2(NET_82),.T3I3(NET_83_CAND3_TRSBL_18_tpGCLKBUF),.TB3S(NET_627),.C3Z(NET_625),.Q3Z(tcdm_result_p2[12]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_R14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_48),.B0I1(m0_m1_dataout_int[31]),.B0I2(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.B0I3(tcdm_result_p2[31]),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[16]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.B0Z(NET_603),.Q0Z(tcdm_result_p2[16]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[31]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R14_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(NET_48),.T2I1(m0_m1_dataout_int[20]),.T2I2(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.T2I3(tcdm_result_p2[20]),.TB2S(GND),.C2Z(NET_386),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_R14_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[20]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T3I0(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.T3I1(tcdm_result_p2[16]),.T3I2(m0_m1_dataout_int[16]),.T3I3(NET_48),.TB3S(GND),.C3Z(NET_312),.Q3Z(tcdm_result_p2[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_R15_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[27]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p2[30]),.T0I1(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.T0I2(NET_48),.T0I3(m0_m1_dataout_int[30]),.TB0S(GND),.C0Z(NET_585),.Q0Z(tcdm_result_p2[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R15_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(NET_19),.T1I1(lint_ADDR_int[7]),.T1I2(NET_15),.T1I3(lint_ADDR_int[2]),.C1Z(NET_52),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_R15_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.B2I1(tcdm_result_p2[25]),.B2I2(NET_48),.B2I3(m0_m1_dataout_int[25]),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.T2I1(m0_m1_dataout_int[27]),.T2I2(NET_48),.T2I3(tcdm_result_p2[27]),.TB2S(GND),.B2Z(NET_496),.C2Z(NET_532),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_R15_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[25]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T3I0(NET_7),.T3I1(NET_14),.T3I2(GND),.T3I3(GND),.C3Z(NET_48),.Q3Z(tcdm_result_p2[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_R16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R16_1 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(NET_15),.T1I2(NET_10),.T1I3(GND),.C1Z(NET_35),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_R16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R16_3 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[30]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(GND),.T3I2(NET_10),.T3I3(NET_7),.TB3S(GND),.C3Z(NET_34),.Q3Z(tcdm_result_p2[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_S11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S11_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_m1_dataout_int[23]),.T1I1(m1_m1_dataout_int[23]),.T1I2(NET_86),.T1I3(NET_83_CAND3_TRSBL_19_tpGCLKBUF),.TB1S(GND),.C1Z(NET_443),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_S11_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_83_CAND3_TRSBL_19_tpGCLKBUF),.T2I1(m1_m1_dataout_int[19]),.T2I2(NET_86),.T2I3(m0_m1_dataout_int[19]),.TB2S(GND),.C2Z(NET_372),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S12_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_83_CAND3_TRSBL_19_tpGCLKBUF),.B0I1(m1_m1_dataout_int[22]),.B0I2(NET_86),.B0I3(m0_m1_dataout_int[22]),.T0I0(m0_m1_dataout_int[18]),.T0I1(NET_86),.T0I2(NET_83_CAND3_TRSBL_19_tpGCLKBUF),.T0I3(m1_m1_dataout_int[18]),.TB0S(GND),.B0Z(NET_425),.C0Z(NET_353),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_S12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S12_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_83_CAND3_TRSBL_19_tpGCLKBUF),.B2I1(NET_86),.B2I2(m1_m1_dataout_int[17]),.B2I3(m0_m1_dataout_int[17]),.T2I0(m0_m1_dataout_int[21]),.T2I1(m1_m1_dataout_int[21]),.T2I2(NET_83_CAND3_TRSBL_19_tpGCLKBUF),.T2I3(NET_86),.TB2S(GND),.B2Z(NET_335),.C2Z(NET_407),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S13_0 (.tFragBitInfo(16'b0101111100000000),.bFragBitInfo(16'b0001001100000000),.B0I0(NET_52_CAND2_TRSBL_19_tpGCLKBUF),.B0I1(tcdm_result_p1[14]),.B0I2(m0_m1_dataout_int[14]),.B0I3(NET_736),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[14]),.Q0EN(tcdm_valid_p1_int_CAND5_TRSBL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T0I0(NET_52_CAND2_TRSBL_19_tpGCLKBUF),.T0I1(tcdm_result_p1[14]),.T0I2(m0_m1_dataout_int[14]),.T0I3(NET_736),.TB0S(NET_50_CAND4_TRSBL_19_tpGCLKBUF),.C0Z(NET_737),.Q0Z(tcdm_result_p1[14]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S13_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[2]),.T1I1(lint_ADDR_int[7]),.T1I2(NET_87),.T1I3(NET_7),.TB1S(GND),.C1Z(NET_83),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_S13_2 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0000000000101010),.B2I0(NET_740),.B2I1(m0_m1_dataout_int[15]),.B2I2(NET_52_CAND2_TRSBL_19_tpGCLKBUF),.B2I3(tcdm_result_p1[15]),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[15]),.Q2EN(tcdm_valid_p1_int_CAND5_TRSBL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T2I0(NET_740),.T2I1(m0_m1_dataout_int[15]),.T2I2(NET_52_CAND2_TRSBL_19_tpGCLKBUF),.T2I3(tcdm_result_p1[15]),.TB2S(NET_50_CAND4_TRSBL_19_tpGCLKBUF),.C2Z(NET_741),.Q2Z(tcdm_result_p1[15]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_S13_3 (.tFragBitInfo(16'b0111011100000000),.bFragBitInfo(16'b0000010001000100),.B3I0(tcdm_result_p1[11]),.B3I1(NET_732),.B3I2(NET_52_CAND2_TRSBL_19_tpGCLKBUF),.B3I3(m0_m1_dataout_int[11]),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[11]),.Q3EN(tcdm_valid_p1_int_CAND5_TRSBL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T3I0(NET_52_CAND2_TRSBL_19_tpGCLKBUF),.T3I1(m0_m1_dataout_int[11]),.T3I2(tcdm_result_p1[11]),.T3I3(NET_732),.TB3S(NET_50_CAND4_TRSBL_19_tpGCLKBUF),.C3Z(NET_733),.Q3Z(tcdm_result_p1[11]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_S16_0 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0001111101011111),.B0I0(tcdm_result_p2[11]),.B0I1(NET_49),.B0I2(NET_7),.B0I3(tcdm_result_p3[11]),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p2[11]),.T0I1(NET_49),.T0I2(NET_7),.T0I3(tcdm_result_p3[11]),.TB0S(NET_14),.C0Z(NET_732),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S16_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[11]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T1I0(NET_35),.T1I1(tcdm_rdata_p1_int[11]),.T1I2(tcdm_rdata_p3_int[11]),.T1I3(NET_34),.TB1S(GND),.C1Z(NET_200),.Q1Z(tcdm_result_p3[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_S16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[11]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p2[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_S16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S17_0 (.tFragBitInfo(16'b0111011111111111),.bFragBitInfo(16'b0000011111111111),.B0I0(NET_49_CAND2_BRSTL_19_tpGCLKBUF),.B0I1(tcdm_result_p3[15]),.B0I2(tcdm_result_p2[15]),.B0I3(NET_7_CAND3_BRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.T0I0(NET_49_CAND2_BRSTL_19_tpGCLKBUF),.T0I1(tcdm_result_p3[15]),.T0I2(tcdm_result_p2[15]),.T0I3(NET_7_CAND3_BRSTL_19_tpGCLKBUF),.TB0S(NET_14),.C0Z(NET_740),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[15]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S17_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B2I0(tcdm_rdata_p1_int[14]),.B2I1(tcdm_rdata_p3_int[14]),.B2I2(NET_34),.B2I3(NET_35),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[15]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(NET_35),.T2I1(tcdm_rdata_p3_int[15]),.T2I2(NET_34),.T2I3(tcdm_rdata_p1_int[15]),.TB2S(GND),.B2Z(NET_260),.C2Z(NET_298),.Q2Z(tcdm_result_p3[15]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_S17_3 (.tFragBitInfo(16'b0101111111111111),.bFragBitInfo(16'b0011001101111111),.B3I0(tcdm_result_p3[14]),.B3I1(NET_7_CAND3_BRSTL_19_tpGCLKBUF),.B3I2(NET_49_CAND2_BRSTL_19_tpGCLKBUF),.B3I3(tcdm_result_p2[14]),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[14]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.T3I0(NET_49_CAND2_BRSTL_19_tpGCLKBUF),.T3I1(tcdm_result_p2[14]),.T3I2(tcdm_result_p3[14]),.T3I3(NET_7_CAND3_BRSTL_19_tpGCLKBUF),.TB3S(NET_14),.C3Z(NET_736),.Q3Z(tcdm_result_p3[14]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_S18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[14]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_S18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_T12_0 (.tFragBitInfo(16'b0101000011110000),.bFragBitInfo(16'b0001000000110000),.B0I0(m0_m1_dataout_int[5]),.B0I1(tcdm_result_p1[5]),.B0I2(NET_756),.B0I3(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[5]),.Q0EN(tcdm_valid_p1_int_CAND5_TRSBL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T0I0(m0_m1_dataout_int[5]),.T0I1(tcdm_result_p1[5]),.T0I2(NET_756),.T0I3(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.TB0S(NET_50_CAND4_TRSBL_20_tpGCLKBUF),.C0Z(NET_757),.Q0Z(tcdm_result_p1[5]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[13]),.Q1EN(tcdm_valid_p1_int_CAND5_TRSBL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p1[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_T12_3 (.tFragBitInfo(16'b0100010011001100),.bFragBitInfo(16'b0001010100000000),.B3I0(tcdm_result_p1[13]),.B3I1(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.B3I2(m0_m1_dataout_int[13]),.B3I3(NET_734),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T3I0(m0_m1_dataout_int[13]),.T3I1(NET_734),.T3I2(tcdm_result_p1[13]),.T3I3(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.TB3S(NET_50_CAND4_TRSBL_20_tpGCLKBUF),.C3Z(NET_735),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_T14_0 (.tFragBitInfo(16'b0100110001001100),.bFragBitInfo(16'b0000000001001100),.B0I0(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.B0I1(NET_728),.B0I2(m0_m1_dataout_int[9]),.B0I3(tcdm_result_p1[9]),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T0I0(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.T0I1(NET_728),.T0I2(m0_m1_dataout_int[9]),.T0I3(tcdm_result_p1[9]),.TB0S(NET_50_CAND4_TRSBL_20_tpGCLKBUF),.C0Z(NET_729),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_T14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[9]),.Q3EN(tcdm_valid_p1_int_CAND5_TRSBL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p1[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_T16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[5]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p3[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T16_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p3_int[5]),.T1I1(tcdm_rdata_p1_int[5]),.T1I2(NET_35),.T1I3(NET_34),.TB1S(GND),.C1Z(NET_653),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_T16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_T16_3 (.tFragBitInfo(16'b0111011111111111),.bFragBitInfo(16'b0001111101011111),.B3I0(tcdm_result_p2[5]),.B3I1(tcdm_result_p3[5]),.B3I2(NET_7),.B3I3(NET_49),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T3I0(NET_7),.T3I1(NET_49),.T3I2(tcdm_result_p2[5]),.T3I3(tcdm_result_p3[5]),.TB3S(NET_14),.C3Z(NET_756),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_T17_0 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0011011101110111),.B0I0(tcdm_result_p2[13]),.B0I1(NET_7_CAND3_BRSTL_20_tpGCLKBUF),.B0I2(NET_49_CAND2_BRSTL_20_tpGCLKBUF),.B0I3(tcdm_result_p3[13]),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[9]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p2[13]),.T0I1(NET_7_CAND3_BRSTL_20_tpGCLKBUF),.T0I2(NET_49_CAND2_BRSTL_20_tpGCLKBUF),.T0I3(tcdm_result_p3[13]),.TB0S(NET_14),.C0Z(NET_734),.Q0Z(tcdm_result_p3[9]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T17_1 (.tFragBitInfo(16'b0111111101111111),.bFragBitInfo(16'b0001001111111111),.B1I0(NET_49_CAND2_BRSTL_20_tpGCLKBUF),.B1I1(tcdm_result_p2[9]),.B1I2(tcdm_result_p3[9]),.B1I3(NET_7_CAND3_BRSTL_20_tpGCLKBUF),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[13]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p3[9]),.T1I1(NET_7_CAND3_BRSTL_20_tpGCLKBUF),.T1I2(NET_49_CAND2_BRSTL_20_tpGCLKBUF),.T1I3(tcdm_result_p2[9]),.TB1S(NET_14),.C1Z(NET_728),.Q1Z(tcdm_result_p3[13]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_T17_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000010000000000),.B2I0(GND),.B2I1(lint_ADDR_int[2]),.B2I2(GND),.B2I3(lint_ADDR_int[3]),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p1_int[9]),.T2I1(tcdm_rdata_p3_int[9]),.T2I2(NET_34),.T2I3(NET_35),.TB2S(GND),.B2Z(NET_131),.C2Z(NET_158),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_T17_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[5]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p3_int[13]),.T3I1(NET_34),.T3I2(tcdm_rdata_p1_int[13]),.T3I3(NET_35),.TB3S(GND),.C3Z(NET_240),.Q3Z(tcdm_result_p2[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_T18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[9]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p2[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[13]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_T18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_U12_0 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0000000000101010),.B0I0(NET_760),.B0I1(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.B0I2(m0_m1_dataout_int[3]),.B0I3(tcdm_result_p1[3]),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[4]),.Q0EN(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T0I0(NET_760),.T0I1(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.T0I2(m0_m1_dataout_int[3]),.T0I3(tcdm_result_p1[3]),.TB0S(NET_50_CAND4_TRSBL_21_tpGCLKBUF),.C0Z(NET_761),.Q0Z(tcdm_result_p1[4]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[3]),.Q1EN(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p1[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U12_2 (.tFragBitInfo(16'b0000101010101010),.bFragBitInfo(16'b0000001000100010),.B2I0(NET_758),.B2I1(tcdm_result_p1[4]),.B2I2(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.B2I3(m0_m1_dataout_int[4]),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[1]),.Q2EN(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T2I0(NET_758),.T2I1(tcdm_result_p1[4]),.T2I2(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.T2I3(m0_m1_dataout_int[4]),.TB2S(NET_50_CAND4_TRSBL_21_tpGCLKBUF),.C2Z(NET_759),.Q2Z(tcdm_result_p1[1]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_U12_3 (.tFragBitInfo(16'b0011000011110000),.bFragBitInfo(16'b0000001000001010),.B3I0(NET_726),.B3I1(m0_m1_dataout_int[1]),.B3I2(tcdm_result_p1[1]),.B3I3(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p1[1]),.T3I1(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.T3I2(NET_726),.T3I3(m0_m1_dataout_int[1]),.TB3S(NET_50_CAND4_TRSBL_21_tpGCLKBUF),.C3Z(NET_727),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_U13_0 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[4]),.T0I1(lint_ADDR_int[5]),.T0I2(lint_ADDR_int[3]),.T0I3(lint_ADDR_int[6]),.TB0S(GND),.C0Z(NET_7),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[10]),.Q2EN(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p1[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U13_3 (.tFragBitInfo(16'b0000101010101010),.bFragBitInfo(16'b0000000001110000),.B3I0(m0_m1_dataout_int[10]),.B3I1(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.B3I2(NET_730),.B3I3(tcdm_result_p1[10]),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(NET_730),.T3I1(tcdm_result_p1[10]),.T3I2(m0_m1_dataout_int[10]),.T3I3(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.TB3S(NET_50_CAND4_TRSBL_21_tpGCLKBUF),.C3Z(NET_731),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_U14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U14_1 (.tFragBitInfo(16'b0010001010101010),.bFragBitInfo(16'b0001000001010000),.B1I0(tcdm_result_p1[8]),.B1I1(m0_m1_dataout_int[8]),.B1I2(NET_738),.B1I3(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[8]),.Q1EN(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T1I0(NET_738),.T1I1(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.T1I2(tcdm_result_p1[8]),.T1I3(m0_m1_dataout_int[8]),.TB1S(NET_50_CAND4_TRSBL_21_tpGCLKBUF),.C1Z(NET_739),.Q1Z(tcdm_result_p1[8]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_U14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_U15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[3]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p2[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U15_3 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0011011100111111),.B3I0(tcdm_result_p3[3]),.B3I1(NET_7),.B3I2(tcdm_result_p2[3]),.B3I3(NET_49),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p2[3]),.T3I1(NET_49),.T3I2(tcdm_result_p3[3]),.T3I3(NET_7),.TB3S(NET_14),.C3Z(NET_760),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_U16_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B0I0(tcdm_rdata_p1_int[4]),.B0I1(NET_34),.B0I2(tcdm_rdata_p3_int[4]),.B0I3(NET_35),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T0I0(NET_34),.T0I1(tcdm_rdata_p3_int[10]),.T0I2(tcdm_rdata_p1_int[10]),.T0I3(NET_35),.TB0S(GND),.B0Z(NET_673),.C0Z(NET_181),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U16_1 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0011011100111111),.B1I0(tcdm_result_p3[4]),.B1I1(NET_7),.B1I2(tcdm_result_p2[4]),.B1I3(NET_49),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[3]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p2[4]),.T1I1(NET_49),.T1I2(tcdm_result_p3[4]),.T1I3(NET_7),.TB1S(NET_14),.C1Z(NET_758),.Q1Z(tcdm_result_p3[3]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_U16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_34),.B2I1(tcdm_rdata_p1_int[1]),.B2I2(tcdm_rdata_p3_int[1]),.B2I3(NET_35),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[4]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B2Z(NET_24),.Q2Z(tcdm_result_p2[4]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U16_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[4]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(NET_34),.T3I1(NET_35),.T3I2(tcdm_rdata_p3_int[3]),.T3I3(tcdm_rdata_p1_int[3]),.C3Z(NET_692),.Q3Z(tcdm_result_p3[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_U17_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[1]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.T0I0(NET_34),.T0I1(tcdm_rdata_p3_int[8]),.T0I2(NET_35),.T0I3(tcdm_rdata_p1_int[8]),.TB0S(GND),.C0Z(NET_279),.Q0Z(tcdm_result_p2[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U17_1 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0101011101011111),.B1I0(NET_7_CAND3_BRSTL_21_tpGCLKBUF),.B1I1(NET_49_CAND2_BRSTL_21_tpGCLKBUF),.B1I2(tcdm_result_p2[10]),.B1I3(tcdm_result_p3[10]),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[8]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p2[10]),.T1I1(tcdm_result_p3[10]),.T1I2(NET_7_CAND3_BRSTL_21_tpGCLKBUF),.T1I3(NET_49_CAND2_BRSTL_21_tpGCLKBUF),.TB1S(NET_14),.C1Z(NET_730),.Q1Z(tcdm_result_p3[8]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_U17_2 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0001111101011111),.B2I0(tcdm_result_p2[1]),.B2I1(NET_49_CAND2_BRSTL_21_tpGCLKBUF),.B2I2(NET_7_CAND3_BRSTL_21_tpGCLKBUF),.B2I3(tcdm_result_p3[1]),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[10]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p2[1]),.T2I1(NET_49_CAND2_BRSTL_21_tpGCLKBUF),.T2I2(NET_7_CAND3_BRSTL_21_tpGCLKBUF),.T2I3(tcdm_result_p3[1]),.TB2S(NET_14),.C2Z(NET_726),.Q2Z(tcdm_result_p3[10]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_U17_3 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0011011100111111),.B3I0(tcdm_result_p3[8]),.B3I1(NET_7_CAND3_BRSTL_21_tpGCLKBUF),.B3I2(tcdm_result_p2[8]),.B3I3(NET_49_CAND2_BRSTL_21_tpGCLKBUF),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[1]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p2[8]),.T3I1(NET_49_CAND2_BRSTL_21_tpGCLKBUF),.T3I2(tcdm_result_p3[8]),.T3I3(NET_7_CAND3_BRSTL_21_tpGCLKBUF),.TB3S(NET_14),.C3Z(NET_738),.Q3Z(tcdm_result_p3[1]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_U18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[8]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p2[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[10]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p2[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V13_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(RESET_int[0]),.TB2S(GND),.C2Z(not_RESET_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_V13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V16_3 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(GND),.T3I1(lint_ADDR_int[3]),.T3I2(NET_65),.T3I3(GND),.C3Z(NET_644),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_W19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(NET_762),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx25587z1),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx25587z1),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx30664z1),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[30]),.Q2EN(nx30664z1),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[30]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[23]),.Q2EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[24]),.Q3EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[19]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[22]),.Q0EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[26]),.Q1EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[13]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[27]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[29]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[21]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[1]),.Q0EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_waddr_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[0]),.Q2EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_waddr_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[3]),.Q0EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_waddr_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[4]),.Q1EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_waddr_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[0]),.Q2EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_waddr_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[7]),.Q3EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_waddr_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[5]),.Q0EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_waddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[8]),.Q1EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_waddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[11]),.Q2EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_waddr_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[11]),.Q3EN(nx18281z1_CAND5_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_raddr_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[6]),.Q0EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_waddr_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[2]),.Q1EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_waddr_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[8]),.Q1EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_waddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[11]),.Q3EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_waddr_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[11]),.Q0EN(nx53672z1_CAND4_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_raddr_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[6]),.Q1EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_waddr_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[2]),.Q2EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_waddr_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[3]),.Q3EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_waddr_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[9]),.Q0EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_waddr_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[7]),.Q1EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_waddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[10]),.Q2EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_waddr_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[4]),.Q3EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_waddr_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[9]),.Q0EN(nx25587z1_CAND2_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_waddr_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[10]),.Q1EN(nx25587z1_CAND2_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_waddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[0]),.Q2EN(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_raddr_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_raddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(NET_762),.Q0EN(nx25587z1_CAND2_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_we_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[8]),.Q2EN(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_raddr_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[6]),.Q3EN(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_raddr_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB11_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(lint_ADDR_int[2]),.T2I1(GND),.T2I2(GND),.T2I3(NET_65),.TB2S(GND),.C2Z(NET_145),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_AB11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[8]),.Q0EN(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_raddr_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[6]),.Q0EN(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_raddr_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(NET_762),.Q2EN(nx30664z1_CAND5_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_we_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[0]),.Q0EN(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_raddr_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[5]),.Q1EN(nx30664z1_CAND5_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_waddr_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[1]),.Q2EN(nx30664z1_CAND5_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_waddr_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_raddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[1]),.Q0EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_raddr_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[3]),.Q1EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_raddr_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[4]),.Q2EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_raddr_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[9]),.Q3EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_raddr_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[7]),.Q1EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_raddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[5]),.Q2EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_raddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[2]),.Q3EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_raddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx41193z1_CAND3_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B0I0(NET_65),.B0I1(lint_ADDR_int[3]),.B0I2(lint_ADDR_int[2]),.B0I3(NET_173),.T0I0(NET_65),.T0I1(lint_ADDR_int[3]),.T0I2(lint_ADDR_int[2]),.T0I3(NET_173),.TB0S(lint_ADDR_int[7]),.C0Z(nx41193z1),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_AC8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC9_0 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b1110101010101010),.B0I0(tcdm_gnt_p1_int),.B0I1(NET_136),.B0I2(NET_133),.B0I3(NET_132),.CD0S(GND),.Q0DI(GND),.Q0EN(nx11312z2),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(NET_136),.T0I2(NET_133),.T0I3(NET_132),.TB0S(GND),.B0Z(nx11312z2),.Q0Z(tcdm_req_p1_dup_0),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AC9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC9_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.T3I0(NET_65),.T3I1(lint_ADDR_int[2]),.T3I2(GND),.T3I3(lint_ADDR_int[3]),.C3Z(NET_136),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_AC10_0 (.tFragBitInfo(16'b0000000000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx36058z1_CAND2_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.T0I0(NET_65),.T0I1(lint_ADDR_int[2]),.T0I2(lint_ADDR_int[3]),.T0I3(GND),.TB0S(GND),.C0Z(NET_137),.Q0Z(tcdm_wdata_p1_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AC10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1111100011110000),.B2I0(NET_132),.B2I1(NET_137),.B2I2(tcdm_gnt_p0_int),.B2I3(NET_133),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx36058z1_CAND2_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B2Z(nx11313z3),.Q2Z(tcdm_wdata_p1_dup_0[6]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC10_3 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx11313z3),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.T3I0(NET_132),.T3I1(NET_137),.T3I2(GND),.T3I3(NET_133),.TB3S(GND),.Q3Z(tcdm_req_p0_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AC12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[23]),.Q2EN(nx36058z1_CAND2_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000010000000),.B0I0(NET_173),.B0I1(NET_65),.B0I2(lint_ADDR_int[2]),.B0I3(lint_ADDR_int[3]),.T0I0(NET_173),.T0I1(NET_65),.T0I2(lint_ADDR_int[2]),.T0I3(lint_ADDR_int[3]),.TB0S(lint_ADDR_int[7]),.C0Z(nx36058z1),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_AC13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC13_3 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int[5]),.T3I1(lint_ADDR_int[4]),.T3I2(lint_ADDR_int[7]),.T3I3(GND),.C3Z(NET_132),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_AC16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001000),.B0I0(RESET_int[0]),.B0I1(NET_65),.B0I2(lint_ADDR_int[5]),.B0I3(lint_ADDR_int[4]),.T0I0(RESET_int[0]),.T0I1(NET_65),.T0I2(lint_ADDR_int[5]),.T0I3(lint_ADDR_int[4]),.TB0S(NET_131),.C0Z(NET_666),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_AC16_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_666),.T1I1(NET_133),.T1I2(NET_147),.T1I3(GND),.TB1S(GND),.C1Z(nx65467z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_AC16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC17_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000001000),.B0I0(lint_ADDR_int[3]),.B0I1(NET_65),.B0I2(lint_ADDR_int[2]),.B0I3(GND),.CD0S(GND),.Q0DI(GND),.Q0EN(nx11310z2),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.T0I0(NET_131),.T0I1(NET_65),.T0I2(NET_133),.T0I3(NET_132),.TB0S(GND),.B0Z(NET_135),.Q0Z(tcdm_req_p3_dup_0),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AC17_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx11311z2),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.T1I0(NET_133),.T1I1(lint_ADDR_int[3]),.T1I2(NET_134),.T1I3(NET_132),.TB1S(GND),.Q1Z(tcdm_req_p2_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AC17_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1110110011001100),.B2I0(NET_133),.B2I1(tcdm_gnt_p2_int),.B2I2(NET_135),.B2I3(NET_132),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.T2I0(NET_131),.T2I1(NET_65),.T2I2(NET_147),.T2I3(NET_173),.TB2S(GND),.B2Z(nx11311z2),.C2Z(nx2520z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_AC17_3 (.tFragBitInfo(16'b1111000011110000),.bFragBitInfo(16'b1110101010101010),.B3I0(tcdm_gnt_p3_int),.B3I1(NET_132),.B3I2(NET_131),.B3I3(NET_65),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.T3I0(NET_131),.T3I1(NET_65),.T3I2(tcdm_gnt_p3_int),.T3I3(NET_132),.TB3S(NET_133),.C3Z(nx11310z2),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_AC18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_131),.B0I1(lint_ADDR_int[7]),.B0I2(NET_65),.B0I3(NET_173),.B0Z(nx25788z1),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000010000000),.B3I0(lint_ADDR_int[3]),.B3I1(NET_173),.B3I2(NET_65),.B3I3(lint_ADDR_int[2]),.T3I0(NET_65),.T3I1(lint_ADDR_int[2]),.T3I2(lint_ADDR_int[3]),.T3I3(NET_173),.TB3S(lint_ADDR_int[7]),.C3Z(nx30923z1),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_AC20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx30923z1_CAND4_BRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[23]),.Q2EN(nx25788z1_CAND3_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[1]),.Q0EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_raddr_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[2]),.Q2EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_raddr_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[3]),.Q3EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_raddr_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[5]),.Q0EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_raddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[7]),.Q1EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_raddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[4]),.Q2EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_raddr_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[9]),.Q3EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_raddr_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx47611z1_CAND4_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[13]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx47611z1_CAND4_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx47611z1_CAND4_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p0_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[20]),.Q2EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[20]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(GND),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(GND),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(GND),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_BE_int[2]),.Q3EN(nx25326z1),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_be_p0_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_BE_int[2]),.Q0EN(nx16907z1),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_be_p1_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx16907z1),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_wen_p1_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD10_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx52746z1_CAND3_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.T1I0(NET_68),.T1I1(RESET_int[0]),.T1I2(NET_174),.T1I3(NET_147),.TB1S(GND),.C1Z(nx25326z1),.Q1Z(tcdm_addr_p1_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_AD10_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx52746z1_CAND3_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.T2I0(NET_145),.T2I1(NET_146),.T2I2(RESET_int[0]),.T2I3(NET_147),.TB2S(GND),.C2Z(nx16907z1),.Q2Z(tcdm_addr_p1_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_AD10_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.T3I0(NET_68),.T3I1(GND),.T3I2(NET_174),.T3I3(NET_147),.TB3S(GND),.C3Z(nx47611z1),.Q3Z(tcdm_wdata_p1_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_AD11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx52746z1_CAND3_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p1_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[21]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD12_3 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx52746z1_CAND3_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_147),.T3I2(NET_145),.T3I3(NET_146),.TB3S(GND),.C3Z(nx52746z1),.Q3Z(tcdm_addr_p1_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_AD13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000000000000),.B0I0(NET_147),.B0I1(GND),.B0I2(NET_68),.B0I3(NET_644),.B0Z(nx57881z1),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD16_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_147),.T1I1(RESET_int[0]),.T1I2(NET_68),.T1I3(NET_644),.C1Z(nx8488z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_AD16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_BE_int[2]),.Q1EN(nx8488z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_be_p2_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_BE_int[2]),.Q3EN(nx65467z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_be_p3_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx57881z1_CAND3_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p2_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx57881z1_CAND3_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[13]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx57881z1_CAND3_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx57881z1_CAND3_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p2_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[20]),.Q3EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx2520z1_CAND2_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p3_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx2520z1_CAND2_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p3_dup_0[12]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p3_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx2520z1_CAND2_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p3_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[22]),.Q0EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p3_dup_0[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[21]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p0_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p0_dup_0[19]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx25326z1),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_wen_p0_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(GND),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_BE_int[3]),.Q2EN(nx25326z1),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_be_p0_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_BE_int[1]),.Q3EN(nx25326z1),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_be_p0_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_BE_int[3]),.Q0EN(nx16907z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_be_p1_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_BE_int[0]),.Q1EN(nx25326z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_be_p0_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_BE_int[1]),.Q2EN(nx16907z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_be_p1_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_BE_int[0]),.Q3EN(nx16907z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_be_p1_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p1_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p1_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p1_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[19]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[18]),.Q2EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[18]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p1_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[26]),.Q1EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_BE_int[1]),.Q0EN(nx8488z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_be_p2_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_BE_int[1]),.Q1EN(nx65467z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_be_p3_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_BE_int[3]),.Q2EN(nx8488z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_be_p2_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_BE_int[3]),.Q3EN(nx65467z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_be_p3_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx65467z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_wen_p3_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx8488z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_wen_p2_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_BE_int[0]),.Q2EN(nx8488z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_be_p2_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_BE_int[0]),.Q3EN(nx65467z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_be_p3_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p2_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p2_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p2_dup_0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p2_dup_0[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx2520z1_CAND2_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p3_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx2520z1_CAND2_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[13]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[19]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p3_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p3_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p3_dup_0[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p0_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p0_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p0_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p1_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p1_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p1_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p1_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p1_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p1_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p1_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p1_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[31]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx57881z1),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx57881z1),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p2_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p2_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p2_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p2_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p2_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[8]),.Q1EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[17]),.Q0EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p2_dup_0[17]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p2_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p2_dup_0[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[31]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p3_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p3_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p3_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p3_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p3_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx2520z1_CAND2_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p3_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p3_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx2520z1_CAND2_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p3_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx2520z1_CAND2_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx2520z1_CAND2_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p3_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[25]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p3_dup_0[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	CLOCK QL_INST_IO_CLK0 (.CEN(VCC),.IP(CLK[0]),.IC(CLK_int[0]),.OP());

	CLOCK QL_INST_IO_CLK1 (.CEN(VCC),.IP(CLK[1]),.IC(CLK_int[1]),.OP());

	CLOCK QL_INST_IO_CLK2 (.CEN(VCC),.IP(CLK[2]),.IC(CLK_int[2]),.OP());

	CLOCK QL_INST_IO_CLK3 (.CEN(VCC),.IP(CLK[3]),.IC(CLK_int[3]),.OP());

	CLOCK QL_INST_IO_CLK4 (.CEN(VCC),.IP(CLK[4]),.IC(CLK_int[4]),.OP());

	CLOCK QL_INST_IO_CLK5 (.CEN(VCC),.IP(CLK[5]),.IC(CLK_int[5]),.OP());

	GMUX QL_INST_GMUX_0 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[0]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_0__GMUX_0_padClk));

	GMUX QL_INST_GMUX_1 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[1]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_1__GMUX_1_padClk));

	GMUX QL_INST_GMUX_2 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[2]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_2__GMUX_2_padClk));

	GMUX QL_INST_GMUX_3 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[3]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_3__GMUX_3_padClk));

	GMUX QL_INST_GMUX_4 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[4]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_4__GMUX_4_padClk));

	GMUX QL_INST_GMUX_5 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[5]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_5__GMUX_5_padClk));

	QPMUX QL_INST_QMUX_TL0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_TL0_padClk));

	QPMUX QL_INST_QMUX_TL1 (.GMUXIN(CLK_int_1__GMUX_1_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_1__QMUX_TL1_padClk));

	QPMUX QL_INST_QMUX_TL2 (.GMUXIN(CLK_int_2__GMUX_2_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_2__QMUX_TL2_padClk));

	QMUX QL_INST_QMUX_TL3 (.GMUXIN(CLK_int_3__GMUX_3_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_3__QMUX_TL3_padClk));

	QMUX QL_INST_QMUX_TL4 (.GMUXIN(CLK_int_4__GMUX_4_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_4__QMUX_TL4_padClk));

	QMUX QL_INST_QMUX_TL5 (.GMUXIN(CLK_int_5__GMUX_5_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_5__QMUX_TL5_padClk));

	QPMUX QL_INST_QMUX_TR0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_TR0_padClk));

	QPMUX QL_INST_QMUX_TR1 (.GMUXIN(GND),.IS0(VCC),.IS1(VCC),.QCLKIN(GND),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_TR1_tpGCLKBUF));

	QMUX QL_INST_QMUX_BL0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_BL0_padClk));

	QMUX QL_INST_QMUX_BL1 (.GMUXIN(GND),.IS(VCC),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_BL1_tpGCLKBUF));

	QMUX QL_INST_QMUX_BL2 (.GMUXIN(GND),.IS(VCC),.QHSCK(nx9707z1),.IZ(nx9707z1_QMUX_BL2_tpGCLKBUF));

	QMUX QL_INST_QMUX_BR0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_BR0_padClk));

	QMUX QL_INST_QMUX_BR1 (.GMUXIN(GND),.IS(VCC),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_BR1_tpGCLKBUF));

	QMUX QL_INST_QMUX_BR2 (.GMUXIN(GND),.IS(VCC),.QHSCK(nx2520z1),.IZ(nx2520z1_QMUX_BR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSTL0_padClk));

	SQEMUX QL_INST_SQMUX_TLSTL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(not_RESET_0),.IZ(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx34006z1),.IZ(nx34006z1_SQMUX_TLSTL2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTL3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx44608z1),.IZ(nx44608z1_SQMUX_TLSTL3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTL4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx39840z1),.IZ(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTL5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(lint_ADDR_int[11]),.IZ(lint_ADDR_int_11__SQMUX_TLSTL5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSTR0_padClk));

	SQEMUX QL_INST_SQMUX_TLSTR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(not_RESET_0),.IZ(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx15998z1),.IZ(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTR3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_46),.IZ(NET_46_SQMUX_TLSTR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTR4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_41),.IZ(NET_41_SQMUX_TLSTR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTR5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_45),.IZ(NET_45_SQMUX_TLSTR5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSBL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSBL0_padClk));

	SQEMUX QL_INST_SQMUX_TLSBL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_1__QMUX_TL1_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_1__SQMUX_TLSBL1_padClk));

	SQEMUX QL_INST_SQMUX_TLSBL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(not_RESET_0),.IZ(not_RESET_0_SQMUX_TLSBL2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBL3 (.QMUXIN(CLK_int_3__QMUX_TL3_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_3__SQMUX_TLSBL3_padClk));

	SQMUX QL_INST_SQMUX_TLSBL4 (.QMUXIN(CLK_int_4__QMUX_TL4_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_4__SQMUX_TLSBL4_padClk));

	SQMUX QL_INST_SQMUX_TLSBL5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_8),.IZ(NET_8_SQMUX_TLSBL5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSBR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSBR0_padClk));

	SQEMUX QL_INST_SQMUX_TLSBR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(not_RESET_0),.IZ(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSBR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_2__QMUX_TL2_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_2__SQMUX_TLSBR2_padClk));

	SQMUX QL_INST_SQMUX_TLSBR3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_110),.IZ(NET_110_SQMUX_TLSBR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBR4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_125),.IZ(NET_125_SQMUX_TLSBR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBR5 (.QMUXIN(CLK_int_5__QMUX_TL5_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_5__SQMUX_TLSBR5_padClk));

	SQEMUX QL_INST_SQMUX_TRSTL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSTL0_padClk));

	SQEMUX QL_INST_SQMUX_TRSTR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSTR0_padClk));

	SQEMUX QL_INST_SQMUX_TRSTR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSTR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx25587z1),.IZ(nx25587z1_SQMUX_TRSTR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTR3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx41193z1),.IZ(nx41193z1_SQMUX_TRSTR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTR4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx47611z1),.IZ(nx47611z1_SQMUX_TRSTR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTR5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx18281z1),.IZ(nx18281z1_SQMUX_TRSTR5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSBL0_padClk));

	SQEMUX QL_INST_SQMUX_TRSBL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_52),.IZ(NET_52_SQMUX_TRSBL2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBL3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_83),.IZ(NET_83_SQMUX_TRSBL3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBL4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_50),.IZ(NET_50_SQMUX_TRSBL4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBL5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(tcdm_valid_p1_int),.IZ(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSBR0_padClk));

	SQEMUX QL_INST_SQMUX_TRSBR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx36058z1),.IZ(nx36058z1_SQMUX_TRSBR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBR3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx52746z1),.IZ(nx52746z1_SQMUX_TRSBR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTL0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSTL0_padClk));

	SQMUX QL_INST_SQMUX_BLSTL1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTL2 (.QMUXIN(nx9707z1_QMUX_BL2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTL3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_94),.IZ(NET_94_SQMUX_BLSTL3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTL4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_29),.IZ(NET_29_SQMUX_BLSTL4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTL5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx4939z1),.IZ(nx4939z1_SQMUX_BLSTL5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTR0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSTR0_padClk));

	SQMUX QL_INST_SQMUX_BLSTR1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTR2 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_17),.IZ(NET_17_SQMUX_BLSTR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx49871z1),.IZ(nx49871z1_SQMUX_BLSTR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_18),.IZ(NET_18_SQMUX_BLSTR4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTR5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_28),.IZ(NET_28_SQMUX_BLSTR5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBL0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSBL0_padClk));

	SQMUX QL_INST_SQMUX_BLSBL1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBL2 (.QMUXIN(nx9707z1_QMUX_BL2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBL3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx22245z1),.IZ(nx22245z1_SQMUX_BLSBL3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBL4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx60831z1),.IZ(nx60831z1_SQMUX_BLSBL4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBR0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSBR0_padClk));

	SQMUX QL_INST_SQMUX_BLSBR1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBR2 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx33579z1),.IZ(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_43),.IZ(NET_43_SQMUX_BLSBR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_44),.IZ(NET_44_SQMUX_BLSBR4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBR5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_45),.IZ(NET_45_SQMUX_BLSBR5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTL0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSTL0_padClk));

	SQMUX QL_INST_SQMUX_BRSTL1 (.QMUXIN(not_RESET_0_QMUX_BR1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTL2 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_49),.IZ(NET_49_SQMUX_BRSTL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTL3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_7),.IZ(NET_7_SQMUX_BRSTL3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTR0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSTR0_padClk));

	SQMUX QL_INST_SQMUX_BRSTR1 (.QMUXIN(not_RESET_0_QMUX_BR1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTR2 (.QMUXIN(nx2520z1_QMUX_BR2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(nx2520z1_SQMUX_BRSTR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx57881z1),.IZ(nx57881z1_SQMUX_BRSTR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx30923z1),.IZ(nx30923z1_SQMUX_BRSTR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSBL0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSBL0_padClk));

	SQMUX QL_INST_SQMUX_BRSBR0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSBR0_padClk));

	SQMUX QL_INST_SQMUX_BRSBR1 (.QMUXIN(not_RESET_0_QMUX_BR1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSBR2 (.QMUXIN(nx2520z1_QMUX_BR2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(nx2520z1_SQMUX_BRSBR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx25788z1),.IZ(nx25788z1_SQMUX_BRSBR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx53672z1),.IZ(nx53672z1_SQMUX_BRSBR4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBR5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx30664z1),.IZ(nx30664z1_SQMUX_BRSBR5_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSTL_1 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_1_padClk));

	CAND QL_INST_CAND0_TLSTL_2 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_2_padClk));

	CAND QL_INST_CAND0_TLSTL_3 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_3_padClk));

	CAND QL_INST_CAND0_TLSTL_4 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_4_padClk));

	CAND QL_INST_CAND0_TLSTL_5 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_5_padClk));

	CAND QL_INST_CAND0_TLSTL_6 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_6_padClk));

	CAND QL_INST_CAND0_TLSTL_7 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_7_padClk));

	CAND QL_INST_CAND1_TLSTL_1 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_2 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_3 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_4 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_5 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_6 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_7 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_2 (.CLKIN(nx34006z1_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z1_CAND2_TLSTL_2_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_3 (.CLKIN(nx34006z1_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z1_CAND2_TLSTL_3_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_4 (.CLKIN(nx34006z1_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z1_CAND2_TLSTL_4_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_5 (.CLKIN(nx34006z1_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z1_CAND2_TLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_6 (.CLKIN(nx34006z1_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z1_CAND2_TLSTL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_1 (.CLKIN(nx44608z1_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx44608z1_CAND3_TLSTL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_2 (.CLKIN(nx44608z1_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx44608z1_CAND3_TLSTL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_3 (.CLKIN(nx44608z1_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx44608z1_CAND3_TLSTL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_4 (.CLKIN(nx44608z1_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx44608z1_CAND3_TLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_5 (.CLKIN(nx44608z1_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx44608z1_CAND3_TLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_6 (.CLKIN(nx44608z1_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx44608z1_CAND3_TLSTL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_3 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_4 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_5 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_6 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_7 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTL_4 (.CLKIN(lint_ADDR_int_11__SQMUX_TLSTL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_11__CAND5_TLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTL_5 (.CLKIN(lint_ADDR_int_11__SQMUX_TLSTL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_11__CAND5_TLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTL_8 (.CLKIN(lint_ADDR_int_11__SQMUX_TLSTL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_11__CAND5_TLSTL_8_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSTR_10 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_10_padClk));

	CAND QL_INST_CAND0_TLSTR_11 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_11_padClk));

	CAND QL_INST_CAND0_TLSTR_12 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_12_padClk));

	CAND QL_INST_CAND0_TLSTR_13 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_13_padClk));

	CAND QL_INST_CAND0_TLSTR_14 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_14_padClk));

	CAND QL_INST_CAND0_TLSTR_15 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_15_padClk));

	CAND QL_INST_CAND0_TLSTR_16 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_16_padClk));

	CAND QL_INST_CAND1_TLSTR_10 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_11 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_12 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_13 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_14 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_15 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_16 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_11 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_12 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_13 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_14 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_9 (.CLKIN(NET_46_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_46_CAND3_TLSTR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_10 (.CLKIN(NET_46_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_46_CAND3_TLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_11 (.CLKIN(NET_46_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_46_CAND3_TLSTR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_13 (.CLKIN(NET_46_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_46_CAND3_TLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_14 (.CLKIN(NET_46_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_46_CAND3_TLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_15 (.CLKIN(NET_46_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_46_CAND3_TLSTR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_16 (.CLKIN(NET_46_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_46_CAND3_TLSTR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_10 (.CLKIN(NET_41_SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_41_CAND4_TLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_11 (.CLKIN(NET_41_SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_41_CAND4_TLSTR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_13 (.CLKIN(NET_41_SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_41_CAND4_TLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_14 (.CLKIN(NET_41_SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_41_CAND4_TLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_15 (.CLKIN(NET_41_SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_41_CAND4_TLSTR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_16 (.CLKIN(NET_41_SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_41_CAND4_TLSTR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTR_9 (.CLKIN(NET_45_SQMUX_TLSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_45_CAND5_TLSTR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTR_10 (.CLKIN(NET_45_SQMUX_TLSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_45_CAND5_TLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTR_11 (.CLKIN(NET_45_SQMUX_TLSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_45_CAND5_TLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSBL_0 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_0_padClk));

	CAND QL_INST_CAND0_TLSBL_1 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_1_padClk));

	CAND QL_INST_CAND0_TLSBL_3 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_3_padClk));

	CAND QL_INST_CAND0_TLSBL_4 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_4_padClk));

	CAND QL_INST_CAND0_TLSBL_5 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_5_padClk));

	CAND QL_INST_CAND0_TLSBL_6 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_6_padClk));

	CAND QL_INST_CAND0_TLSBL_7 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_7_padClk));

	CAND QL_INST_CAND0_TLSBL_8 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_8_padClk));

	CAND QL_INST_CAND1_TLSBL_8 (.CLKIN(CLK_int_1__SQMUX_TLSBL1_padClk),.SEN(VCC),.IZ(CLK_int_1__CAND1_TLSBL_8_padClk));

	CAND QL_INST_CAND2_TLSBL_1 (.CLKIN(not_RESET_0_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND2_TLSBL_1_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_3 (.CLKIN(not_RESET_0_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND2_TLSBL_3_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_4 (.CLKIN(not_RESET_0_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND2_TLSBL_4_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_5 (.CLKIN(not_RESET_0_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND2_TLSBL_5_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_6 (.CLKIN(not_RESET_0_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND2_TLSBL_6_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_7 (.CLKIN(not_RESET_0_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND2_TLSBL_7_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_8 (.CLKIN(not_RESET_0_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND2_TLSBL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_5 (.CLKIN(CLK_int_3__SQMUX_TLSBL3_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_3__CAND3_TLSBL_5_padClk));

	CANDEN QL_INST_CAND4_TLSBL_7 (.CLKIN(CLK_int_4__SQMUX_TLSBL4_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_4__CAND4_TLSBL_7_padClk));

	CANDEN QL_INST_CAND5_TLSBL_1 (.CLKIN(NET_8_SQMUX_TLSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_8_CAND5_TLSBL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBL_2 (.CLKIN(NET_8_SQMUX_TLSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_8_CAND5_TLSBL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBL_3 (.CLKIN(NET_8_SQMUX_TLSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_8_CAND5_TLSBL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBL_4 (.CLKIN(NET_8_SQMUX_TLSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_8_CAND5_TLSBL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBL_7 (.CLKIN(NET_8_SQMUX_TLSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_8_CAND5_TLSBL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBL_8 (.CLKIN(NET_8_SQMUX_TLSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_8_CAND5_TLSBL_8_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSBR_9 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_9_padClk));

	CAND QL_INST_CAND0_TLSBR_10 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_10_padClk));

	CAND QL_INST_CAND0_TLSBR_11 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_11_padClk));

	CAND QL_INST_CAND0_TLSBR_12 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_12_padClk));

	CAND QL_INST_CAND0_TLSBR_13 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_13_padClk));

	CAND QL_INST_CAND0_TLSBR_14 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_14_padClk));

	CAND QL_INST_CAND0_TLSBR_15 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_15_padClk));

	CAND QL_INST_CAND0_TLSBR_16 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_16_padClk));

	CAND QL_INST_CAND1_TLSBR_9 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_10 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_11 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_12 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_13 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_14 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_15 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_16 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_9 (.CLKIN(CLK_int_2__SQMUX_TLSBR2_padClk),.SEN(VCC),.IZ(CLK_int_2__CAND2_TLSBR_9_padClk));

	CANDEN QL_INST_CAND3_TLSBR_13 (.CLKIN(NET_110_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_110_CAND3_TLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_14 (.CLKIN(NET_110_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_110_CAND3_TLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_15 (.CLKIN(NET_110_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_110_CAND3_TLSBR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_16 (.CLKIN(NET_110_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_110_CAND3_TLSBR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_13 (.CLKIN(NET_125_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_125_CAND4_TLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_14 (.CLKIN(NET_125_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_125_CAND4_TLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_15 (.CLKIN(NET_125_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_125_CAND4_TLSBR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_16 (.CLKIN(NET_125_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_125_CAND4_TLSBR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBR_9 (.CLKIN(CLK_int_5__SQMUX_TLSBR5_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_5__CAND5_TLSBR_9_padClk));

	CAND QL_INST_CAND0_TRSTL_17 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_17_padClk));

	CAND QL_INST_CAND0_TRSTL_19 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_19_padClk));

	CAND QL_INST_CAND0_TRSTL_24 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_24_padClk));

	CAND QL_INST_CAND0_TRSTR_25 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_25_padClk));

	CAND QL_INST_CAND0_TRSTR_26 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_26_padClk));

	CAND QL_INST_CAND0_TRSTR_27 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_27_padClk));

	CAND QL_INST_CAND0_TRSTR_28 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_28_padClk));

	CAND QL_INST_CAND0_TRSTR_29 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_29_padClk));

	CAND QL_INST_CAND0_TRSTR_30 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_30_padClk));

	CAND QL_INST_CAND0_TRSTR_31 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_31_padClk));

	CAND QL_INST_CAND0_TRSTR_32 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_32_padClk));

	CAND QL_INST_CAND0_TRSTR_33 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_33_padClk));

	CAND QL_INST_CAND1_TRSTR_25 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_26 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_27 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_28 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_29 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_30 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_31 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_32 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTR_25 (.CLKIN(nx25587z1_SQMUX_TRSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTR_26 (.CLKIN(nx25587z1_SQMUX_TRSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTR_27 (.CLKIN(nx25587z1_SQMUX_TRSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTR_28 (.CLKIN(nx25587z1_SQMUX_TRSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx25587z1_CAND2_TRSTR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_29 (.CLKIN(nx41193z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z1_CAND3_TRSTR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_30 (.CLKIN(nx41193z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_31 (.CLKIN(nx41193z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_32 (.CLKIN(nx41193z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_30 (.CLKIN(nx47611z1_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx47611z1_CAND4_TRSTR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_31 (.CLKIN(nx47611z1_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_32 (.CLKIN(nx47611z1_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSTR_27 (.CLKIN(nx18281z1_SQMUX_TRSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx18281z1_CAND5_TRSTR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSTR_28 (.CLKIN(nx18281z1_SQMUX_TRSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSTR_29 (.CLKIN(nx18281z1_SQMUX_TRSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF));

	CAND QL_INST_CAND0_TRSBL_17 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_17_padClk));

	CAND QL_INST_CAND0_TRSBL_18 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_18_padClk));

	CAND QL_INST_CAND0_TRSBL_19 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_19_padClk));

	CAND QL_INST_CAND0_TRSBL_20 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_20_padClk));

	CAND QL_INST_CAND0_TRSBL_21 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_21_padClk));

	CAND QL_INST_CAND1_TRSBL_17 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_18 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_19 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_20 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_21 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBL_18 (.CLKIN(NET_52_SQMUX_TRSBL2_tpGCLKBUF),.SEN(VCC),.IZ(NET_52_CAND2_TRSBL_18_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBL_19 (.CLKIN(NET_52_SQMUX_TRSBL2_tpGCLKBUF),.SEN(VCC),.IZ(NET_52_CAND2_TRSBL_19_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBL_20 (.CLKIN(NET_52_SQMUX_TRSBL2_tpGCLKBUF),.SEN(VCC),.IZ(NET_52_CAND2_TRSBL_20_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBL_21 (.CLKIN(NET_52_SQMUX_TRSBL2_tpGCLKBUF),.SEN(VCC),.IZ(NET_52_CAND2_TRSBL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBL_18 (.CLKIN(NET_83_SQMUX_TRSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_83_CAND3_TRSBL_18_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBL_19 (.CLKIN(NET_83_SQMUX_TRSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_83_CAND3_TRSBL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBL_17 (.CLKIN(NET_50_SQMUX_TRSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_50_CAND4_TRSBL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBL_19 (.CLKIN(NET_50_SQMUX_TRSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_50_CAND4_TRSBL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBL_20 (.CLKIN(NET_50_SQMUX_TRSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_50_CAND4_TRSBL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBL_21 (.CLKIN(NET_50_SQMUX_TRSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_50_CAND4_TRSBL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBL_17 (.CLKIN(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBL_19 (.CLKIN(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p1_int_CAND5_TRSBL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBL_20 (.CLKIN(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p1_int_CAND5_TRSBL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBL_21 (.CLKIN(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF));

	CAND QL_INST_CAND0_TRSBR_29 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_29_padClk));

	CAND QL_INST_CAND0_TRSBR_30 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_30_padClk));

	CAND QL_INST_CAND0_TRSBR_31 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_31_padClk));

	CAND QL_INST_CAND0_TRSBR_32 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_32_padClk));

	CAND QL_INST_CAND0_TRSBR_33 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_33_padClk));

	CAND QL_INST_CAND1_TRSBR_29 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBR_30 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBR_31 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBR_32 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_29 (.CLKIN(nx36058z1_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx36058z1_CAND2_TRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_30 (.CLKIN(nx36058z1_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_31 (.CLKIN(nx36058z1_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_32 (.CLKIN(nx36058z1_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBR_30 (.CLKIN(nx52746z1_SQMUX_TRSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx52746z1_CAND3_TRSBR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBR_31 (.CLKIN(nx52746z1_SQMUX_TRSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBR_32 (.CLKIN(nx52746z1_SQMUX_TRSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSTL_1 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_1_padClk));

	CANDEN QL_INST_CAND0_BLSTL_2 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_2_padClk));

	CANDEN QL_INST_CAND0_BLSTL_3 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_3_padClk));

	CANDEN QL_INST_CAND0_BLSTL_4 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_4_padClk));

	CANDEN QL_INST_CAND0_BLSTL_5 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_5_padClk));

	CANDEN QL_INST_CAND0_BLSTL_6 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_6_padClk));

	CANDEN QL_INST_CAND0_BLSTL_7 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_7_padClk));

	CANDEN QL_INST_CAND0_BLSTL_8 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_8_padClk));

	CANDEN QL_INST_CAND1_BLSTL_1 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_2 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_3 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_4 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_5 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_6 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_7 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_8 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_1 (.CLKIN(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_2 (.CLKIN(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSTL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_3 (.CLKIN(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSTL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_4 (.CLKIN(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_5 (.CLKIN(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_6 (.CLKIN(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSTL_6_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTL_5 (.CLKIN(NET_94_SQMUX_BLSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_94_CAND3_BLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTL_6 (.CLKIN(NET_94_SQMUX_BLSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_94_CAND3_BLSTL_6_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTL_7 (.CLKIN(NET_94_SQMUX_BLSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_94_CAND3_BLSTL_7_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTL_8 (.CLKIN(NET_94_SQMUX_BLSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_94_CAND3_BLSTL_8_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTL_2 (.CLKIN(NET_29_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(NET_29_CAND4_BLSTL_2_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTL_7 (.CLKIN(NET_29_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(NET_29_CAND4_BLSTL_7_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTL_8 (.CLKIN(NET_29_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(NET_29_CAND4_BLSTL_8_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_4 (.CLKIN(nx4939z1_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND5_BLSTL_4_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_5 (.CLKIN(nx4939z1_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND5_BLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_6 (.CLKIN(nx4939z1_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND5_BLSTL_6_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_7 (.CLKIN(nx4939z1_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND5_BLSTL_7_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_8 (.CLKIN(nx4939z1_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND5_BLSTL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSTR_9 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_9_padClk));

	CANDEN QL_INST_CAND0_BLSTR_10 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_10_padClk));

	CANDEN QL_INST_CAND0_BLSTR_11 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_11_padClk));

	CANDEN QL_INST_CAND0_BLSTR_12 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_12_padClk));

	CANDEN QL_INST_CAND0_BLSTR_13 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_13_padClk));

	CANDEN QL_INST_CAND0_BLSTR_14 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_14_padClk));

	CANDEN QL_INST_CAND0_BLSTR_15 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_15_padClk));

	CANDEN QL_INST_CAND1_BLSTR_9 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_10 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_11 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_12 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_13 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_14 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_15 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_9 (.CLKIN(NET_17_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_17_CAND2_BLSTR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_10 (.CLKIN(NET_17_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_17_CAND2_BLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_11 (.CLKIN(NET_17_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_17_CAND2_BLSTR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_12 (.CLKIN(NET_17_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_17_CAND2_BLSTR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_13 (.CLKIN(NET_17_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_17_CAND2_BLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_14 (.CLKIN(NET_17_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_17_CAND2_BLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_9 (.CLKIN(nx49871z1_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx49871z1_CAND3_BLSTR_9_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_10 (.CLKIN(nx49871z1_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx49871z1_CAND3_BLSTR_10_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_11 (.CLKIN(nx49871z1_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx49871z1_CAND3_BLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_12 (.CLKIN(nx49871z1_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx49871z1_CAND3_BLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_13 (.CLKIN(nx49871z1_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx49871z1_CAND3_BLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_14 (.CLKIN(nx49871z1_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx49871z1_CAND3_BLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_9 (.CLKIN(NET_18_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_18_CAND4_BLSTR_9_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_10 (.CLKIN(NET_18_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_18_CAND4_BLSTR_10_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_11 (.CLKIN(NET_18_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_18_CAND4_BLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_9 (.CLKIN(NET_28_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_28_CAND5_BLSTR_9_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_12 (.CLKIN(NET_28_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_28_CAND5_BLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_13 (.CLKIN(NET_28_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_28_CAND5_BLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_14 (.CLKIN(NET_28_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_28_CAND5_BLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSBL_1 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_1_padClk));

	CANDEN QL_INST_CAND0_BLSBL_2 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_2_padClk));

	CANDEN QL_INST_CAND0_BLSBL_3 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_3_padClk));

	CANDEN QL_INST_CAND0_BLSBL_4 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_4_padClk));

	CANDEN QL_INST_CAND0_BLSBL_5 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_5_padClk));

	CANDEN QL_INST_CAND0_BLSBL_6 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_6_padClk));

	CANDEN QL_INST_CAND0_BLSBL_7 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_7_padClk));

	CANDEN QL_INST_CAND0_BLSBL_8 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_8_padClk));

	CANDEN QL_INST_CAND1_BLSBL_1 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_2 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_3 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_4 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_5 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_6 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_7 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_8 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_1 (.CLKIN(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_2 (.CLKIN(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSBL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_3 (.CLKIN(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSBL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_5 (.CLKIN(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSBL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_6 (.CLKIN(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSBL_6_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBL_2 (.CLKIN(nx22245z1_SQMUX_BLSBL3_tpGCLKBUF),.SEN(VCC),.IZ(nx22245z1_CAND3_BLSBL_2_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBL_3 (.CLKIN(nx22245z1_SQMUX_BLSBL3_tpGCLKBUF),.SEN(VCC),.IZ(nx22245z1_CAND3_BLSBL_3_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBL_4 (.CLKIN(nx22245z1_SQMUX_BLSBL3_tpGCLKBUF),.SEN(VCC),.IZ(nx22245z1_CAND3_BLSBL_4_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBL_5 (.CLKIN(nx22245z1_SQMUX_BLSBL3_tpGCLKBUF),.SEN(VCC),.IZ(nx22245z1_CAND3_BLSBL_5_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBL_6 (.CLKIN(nx22245z1_SQMUX_BLSBL3_tpGCLKBUF),.SEN(VCC),.IZ(nx22245z1_CAND3_BLSBL_6_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBL_5 (.CLKIN(nx60831z1_SQMUX_BLSBL4_tpGCLKBUF),.SEN(VCC),.IZ(nx60831z1_CAND4_BLSBL_5_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBL_6 (.CLKIN(nx60831z1_SQMUX_BLSBL4_tpGCLKBUF),.SEN(VCC),.IZ(nx60831z1_CAND4_BLSBL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSBR_9 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_9_padClk));

	CANDEN QL_INST_CAND0_BLSBR_10 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_10_padClk));

	CANDEN QL_INST_CAND0_BLSBR_11 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_11_padClk));

	CANDEN QL_INST_CAND0_BLSBR_12 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_12_padClk));

	CANDEN QL_INST_CAND0_BLSBR_13 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_13_padClk));

	CANDEN QL_INST_CAND0_BLSBR_14 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_14_padClk));

	CANDEN QL_INST_CAND0_BLSBR_15 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_15_padClk));

	CANDEN QL_INST_CAND0_BLSBR_16 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_16_padClk));

	CANDEN QL_INST_CAND1_BLSBR_9 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_10 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_11 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_12 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_13 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_14 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_15 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_16 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_11 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_12 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_13 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_14 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_9 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_9_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_10 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_10_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_11 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_11_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_12 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_12_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_13 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_13_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_14 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_15 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_15_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBR_10 (.CLKIN(NET_44_SQMUX_BLSBR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_44_CAND4_BLSBR_10_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBR_11 (.CLKIN(NET_44_SQMUX_BLSBR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_44_CAND4_BLSBR_11_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBR_12 (.CLKIN(NET_44_SQMUX_BLSBR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_44_CAND4_BLSBR_12_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBR_13 (.CLKIN(NET_44_SQMUX_BLSBR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_44_CAND4_BLSBR_13_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBR_14 (.CLKIN(NET_44_SQMUX_BLSBR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_44_CAND4_BLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBR_15 (.CLKIN(NET_44_SQMUX_BLSBR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_44_CAND4_BLSBR_15_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSBR_9 (.CLKIN(NET_45_SQMUX_BLSBR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_45_CAND5_BLSBR_9_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSBR_10 (.CLKIN(NET_45_SQMUX_BLSBR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_45_CAND5_BLSBR_10_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSBR_11 (.CLKIN(NET_45_SQMUX_BLSBR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_45_CAND5_BLSBR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSTL_19 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_19_padClk));

	CANDEN QL_INST_CAND0_BRSTL_20 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_20_padClk));

	CANDEN QL_INST_CAND0_BRSTL_21 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_21_padClk));

	CANDEN QL_INST_CAND1_BRSTL_19 (.CLKIN(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTL_20 (.CLKIN(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTL_21 (.CLKIN(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_19 (.CLKIN(NET_49_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_49_CAND2_BRSTL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_20 (.CLKIN(NET_49_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_49_CAND2_BRSTL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_21 (.CLKIN(NET_49_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_49_CAND2_BRSTL_21_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTL_19 (.CLKIN(NET_7_SQMUX_BRSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_7_CAND3_BRSTL_19_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTL_20 (.CLKIN(NET_7_SQMUX_BRSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_7_CAND3_BRSTL_20_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTL_21 (.CLKIN(NET_7_SQMUX_BRSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_7_CAND3_BRSTL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSTR_29 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_29_padClk));

	CANDEN QL_INST_CAND0_BRSTR_30 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_30_padClk));

	CANDEN QL_INST_CAND0_BRSTR_31 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_31_padClk));

	CANDEN QL_INST_CAND0_BRSTR_32 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_32_padClk));

	CANDEN QL_INST_CAND0_BRSTR_33 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_33_padClk));

	CANDEN QL_INST_CAND1_BRSTR_29 (.CLKIN(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTR_30 (.CLKIN(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTR_31 (.CLKIN(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTR_32 (.CLKIN(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_30 (.CLKIN(nx2520z1_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSTR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_31 (.CLKIN(nx2520z1_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSTR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_32 (.CLKIN(nx2520z1_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTR_30 (.CLKIN(nx57881z1_SQMUX_BRSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx57881z1_CAND3_BRSTR_30_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTR_31 (.CLKIN(nx57881z1_SQMUX_BRSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTR_32 (.CLKIN(nx57881z1_SQMUX_BRSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTR_29 (.CLKIN(nx30923z1_SQMUX_BRSTR4_tpGCLKBUF),.SEN(VCC),.IZ(nx30923z1_CAND4_BRSTR_29_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTR_30 (.CLKIN(nx30923z1_SQMUX_BRSTR4_tpGCLKBUF),.SEN(VCC),.IZ(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTR_31 (.CLKIN(nx30923z1_SQMUX_BRSTR4_tpGCLKBUF),.SEN(VCC),.IZ(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTR_32 (.CLKIN(nx30923z1_SQMUX_BRSTR4_tpGCLKBUF),.SEN(VCC),.IZ(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSBL_19 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_19_padClk));

	CANDEN QL_INST_CAND0_BRSBL_24 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_24_padClk));

	CANDEN QL_INST_CAND0_BRSBR_25 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_25_padClk));

	CANDEN QL_INST_CAND0_BRSBR_26 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_26_padClk));

	CANDEN QL_INST_CAND0_BRSBR_27 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_27_padClk));

	CANDEN QL_INST_CAND0_BRSBR_28 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_28_padClk));

	CANDEN QL_INST_CAND0_BRSBR_29 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_29_padClk));

	CANDEN QL_INST_CAND0_BRSBR_30 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_30_padClk));

	CANDEN QL_INST_CAND0_BRSBR_31 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_31_padClk));

	CANDEN QL_INST_CAND0_BRSBR_32 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_32_padClk));

	CANDEN QL_INST_CAND1_BRSBR_25 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_26 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_27 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_28 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_29 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_30 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_31 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_32 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_30 (.CLKIN(nx2520z1_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSBR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_31 (.CLKIN(nx2520z1_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_32 (.CLKIN(nx2520z1_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSBR_32_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_29 (.CLKIN(nx25788z1_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z1_CAND3_BRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_30 (.CLKIN(nx25788z1_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_31 (.CLKIN(nx25788z1_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_32 (.CLKIN(nx25788z1_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBR_27 (.CLKIN(nx53672z1_SQMUX_BRSBR4_tpGCLKBUF),.SEN(VCC),.IZ(nx53672z1_CAND4_BRSBR_27_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBR_28 (.CLKIN(nx53672z1_SQMUX_BRSBR4_tpGCLKBUF),.SEN(VCC),.IZ(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBR_29 (.CLKIN(nx53672z1_SQMUX_BRSBR4_tpGCLKBUF),.SEN(VCC),.IZ(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBR_25 (.CLKIN(nx30664z1_SQMUX_BRSBR5_tpGCLKBUF),.SEN(VCC),.IZ(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBR_26 (.CLKIN(nx30664z1_SQMUX_BRSBR5_tpGCLKBUF),.SEN(VCC),.IZ(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBR_27 (.CLKIN(nx30664z1_SQMUX_BRSBR5_tpGCLKBUF),.SEN(VCC),.IZ(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBR_28 (.CLKIN(nx30664z1_SQMUX_BRSBR5_tpGCLKBUF),.SEN(VCC),.IZ(nx30664z1_CAND5_BRSBR_28_tpGCLKBUF));

	OBUF QL_INST_F2A_T_2_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTL_2_padClk),.OUT_OBUF(m0_oper0_wclk));

	OBUF QL_INST_F2A_T_2_1 (.IN_OBUF(m0_oper0_wmode_dup_0[1]),.OUT_OBUF(m0_oper0_wmode[1]));

	OBUF QL_INST_F2A_T_2_2 (.IN_OBUF(m0_oper0_wmode_dup_0[0]),.OUT_OBUF(m0_oper0_wmode[0]));

	OBUF QL_INST_F2A_T_2_3 (.IN_OBUF(m0_oper0_wdsel_dup_0),.OUT_OBUF(m0_oper0_wdsel));

	OBUF QL_INST_F2A_T_2_4 (.IN_OBUF(m0_oper0_rmode_dup_0[1]),.OUT_OBUF(m0_oper0_rmode[1]));

	OBUF QL_INST_F2A_T_2_5 (.IN_OBUF(m0_oper0_rmode_dup_0[0]),.OUT_OBUF(m0_oper0_rmode[0]));

	OBUF QL_INST_F2A_T_2_6 (.IN_OBUF(m0_oper0_wdata_dup_0[31]),.OUT_OBUF(m0_oper0_wdata[31]));

	OBUF QL_INST_F2A_T_2_7 (.IN_OBUF(m0_oper0_wdata_dup_0[30]),.OUT_OBUF(m0_oper0_wdata[30]));

	OBUF QL_INST_F2A_T_2_8 (.IN_OBUF(m0_oper0_wdata_dup_0[29]),.OUT_OBUF(m0_oper0_wdata[29]));

	OBUF QL_INST_F2A_T_2_9 (.IN_OBUF(m0_oper0_wdata_dup_0[28]),.OUT_OBUF(m0_oper0_wdata[28]));

	OBUF QL_INST_F2A_T_2_10 (.IN_OBUF(m0_oper0_wdata_dup_0[27]),.OUT_OBUF(m0_oper0_wdata[27]));

	OBUF QL_INST_F2A_T_2_11 (.IN_OBUF(m0_oper0_wdata_dup_0[26]),.OUT_OBUF(m0_oper0_wdata[26]));

	OBUF QL_INST_F2A_T_2_12 (.IN_OBUF(m0_oper0_wdata_dup_0[25]),.OUT_OBUF(m0_oper0_wdata[25]));

	OBUF QL_INST_F2A_T_2_13 (.IN_OBUF(m0_oper0_wdata_dup_0[24]),.OUT_OBUF(m0_oper0_wdata[24]));

	OBUF QL_INST_F2A_T_2_14 (.IN_OBUF(m0_oper0_wdata_dup_0[23]),.OUT_OBUF(m0_oper0_wdata[23]));

	OBUF QL_INST_F2A_T_2_15 (.IN_OBUF(m0_oper0_wdata_dup_0[22]),.OUT_OBUF(m0_oper0_wdata[22]));

	OBUF QL_INST_F2A_T_2_16 (.IN_OBUF(m0_oper0_wdata_dup_0[21]),.OUT_OBUF(m0_oper0_wdata[21]));

	OBUF QL_INST_F2A_T_2_17 (.IN_OBUF(m0_oper0_wdata_dup_0[20]),.OUT_OBUF(m0_oper0_wdata[20]));

	IBUF QL_INST_A2F_T_2_0 (.IN_IBUF(m0_oper0_rdata[31]),.OUT_IBUF(m0_oper0_rdata_int[31]));

	IBUF QL_INST_A2F_T_2_1 (.IN_IBUF(m0_oper0_rdata[30]),.OUT_IBUF(m0_oper0_rdata_int[30]));

	IBUF QL_INST_A2F_T_2_2 (.IN_IBUF(m0_oper0_rdata[29]),.OUT_IBUF(m0_oper0_rdata_int[29]));

	IBUF QL_INST_A2F_T_2_3 (.IN_IBUF(m0_oper0_rdata[28]),.OUT_IBUF(m0_oper0_rdata_int[28]));

	OBUF QL_INST_F2A_T_3_0 (.IN_OBUF(m0_oper0_wdata_dup_0[19]),.OUT_OBUF(m0_oper0_wdata[19]));

	OBUF QL_INST_F2A_T_3_1 (.IN_OBUF(m0_oper0_wdata_dup_0[18]),.OUT_OBUF(m0_oper0_wdata[18]));

	OBUF QL_INST_F2A_T_3_2 (.IN_OBUF(m0_oper0_wdata_dup_0[17]),.OUT_OBUF(m0_oper0_wdata[17]));

	OBUF QL_INST_F2A_T_3_3 (.IN_OBUF(m0_oper0_wdata_dup_0[16]),.OUT_OBUF(m0_oper0_wdata[16]));

	OBUF QL_INST_F2A_T_3_4 (.IN_OBUF(m0_oper0_wdata_dup_0[15]),.OUT_OBUF(m0_oper0_wdata[15]));

	OBUF QL_INST_F2A_T_3_5 (.IN_OBUF(m0_oper0_wdata_dup_0[14]),.OUT_OBUF(m0_oper0_wdata[14]));

	OBUF QL_INST_F2A_T_3_6 (.IN_OBUF(m0_oper0_wdata_dup_0[13]),.OUT_OBUF(m0_oper0_wdata[13]));

	OBUF QL_INST_F2A_T_3_7 (.IN_OBUF(m0_oper0_wdata_dup_0[12]),.OUT_OBUF(m0_oper0_wdata[12]));

	OBUF QL_INST_F2A_T_3_8 (.IN_OBUF(m0_oper0_wdata_dup_0[11]),.OUT_OBUF(m0_oper0_wdata[11]));

	OBUF QL_INST_F2A_T_3_9 (.IN_OBUF(m0_oper0_wdata_dup_0[10]),.OUT_OBUF(m0_oper0_wdata[10]));

	OBUF QL_INST_F2A_T_3_10 (.IN_OBUF(m0_oper0_wdata_dup_0[9]),.OUT_OBUF(m0_oper0_wdata[9]));

	OBUF QL_INST_F2A_T_3_11 (.IN_OBUF(m0_oper0_wdata_dup_0[8]),.OUT_OBUF(m0_oper0_wdata[8]));

	IBUF QL_INST_A2F_T_3_0 (.IN_IBUF(m0_oper0_rdata[27]),.OUT_IBUF(m0_oper0_rdata_int[27]));

	IBUF QL_INST_A2F_T_3_1 (.IN_IBUF(m0_oper0_rdata[26]),.OUT_IBUF(m0_oper0_rdata_int[26]));

	IBUF QL_INST_A2F_T_3_2 (.IN_IBUF(m0_oper0_rdata[25]),.OUT_IBUF(m0_oper0_rdata_int[25]));

	IBUF QL_INST_A2F_T_3_3 (.IN_IBUF(m0_oper0_rdata[24]),.OUT_IBUF(m0_oper0_rdata_int[24]));

	IBUF QL_INST_A2F_T_3_4 (.IN_IBUF(m0_oper0_rdata[23]),.OUT_IBUF(m0_oper0_rdata_int[23]));

	IBUF QL_INST_A2F_T_3_5 (.IN_IBUF(m0_oper0_rdata[22]),.OUT_IBUF(m0_oper0_rdata_int[22]));

	OBUF QL_INST_F2A_T_4_0 (.IN_OBUF(m0_oper0_wdata_dup_0[7]),.OUT_OBUF(m0_oper0_wdata[7]));

	OBUF QL_INST_F2A_T_4_1 (.IN_OBUF(m0_oper0_wdata_dup_0[6]),.OUT_OBUF(m0_oper0_wdata[6]));

	OBUF QL_INST_F2A_T_4_2 (.IN_OBUF(m0_oper0_wdata_dup_0[5]),.OUT_OBUF(m0_oper0_wdata[5]));

	OBUF QL_INST_F2A_T_4_3 (.IN_OBUF(m0_oper0_wdata_dup_0[4]),.OUT_OBUF(m0_oper0_wdata[4]));

	OBUF QL_INST_F2A_T_4_4 (.IN_OBUF(m0_oper0_wdata_dup_0[3]),.OUT_OBUF(m0_oper0_wdata[3]));

	OBUF QL_INST_F2A_T_4_5 (.IN_OBUF(m0_oper0_wdata_dup_0[2]),.OUT_OBUF(m0_oper0_wdata[2]));

	OBUF QL_INST_F2A_T_4_6 (.IN_OBUF(m0_oper0_wdata_dup_0[1]),.OUT_OBUF(m0_oper0_wdata[1]));

	OBUF QL_INST_F2A_T_4_7 (.IN_OBUF(m0_oper0_wdata_dup_0[0]),.OUT_OBUF(m0_oper0_wdata[0]));

	OBUF QL_INST_F2A_T_4_8 (.IN_OBUF(m0_oper0_waddr_dup_0[11]),.OUT_OBUF(m0_oper0_waddr[11]));

	OBUF QL_INST_F2A_T_4_9 (.IN_OBUF(m0_oper0_waddr_dup_0[10]),.OUT_OBUF(m0_oper0_waddr[10]));

	OBUF QL_INST_F2A_T_4_10 (.IN_OBUF(m0_oper0_waddr_dup_0[9]),.OUT_OBUF(m0_oper0_waddr[9]));

	OBUF QL_INST_F2A_T_4_11 (.IN_OBUF(m0_oper0_waddr_dup_0[8]),.OUT_OBUF(m0_oper0_waddr[8]));

	OBUF QL_INST_F2A_T_4_12 (.IN_OBUF(m0_oper0_waddr_dup_0[7]),.OUT_OBUF(m0_oper0_waddr[7]));

	OBUF QL_INST_F2A_T_4_13 (.IN_OBUF(m0_oper0_waddr_dup_0[6]),.OUT_OBUF(m0_oper0_waddr[6]));

	OBUF QL_INST_F2A_T_4_14 (.IN_OBUF(m0_oper0_waddr_dup_0[5]),.OUT_OBUF(m0_oper0_waddr[5]));

	OBUF QL_INST_F2A_T_4_15 (.IN_OBUF(m0_oper0_waddr_dup_0[4]),.OUT_OBUF(m0_oper0_waddr[4]));

	OBUF QL_INST_F2A_T_4_16 (.IN_OBUF(m0_oper0_waddr_dup_0[3]),.OUT_OBUF(m0_oper0_waddr[3]));

	OBUF QL_INST_F2A_T_4_17 (.IN_OBUF(m0_oper0_waddr_dup_0[2]),.OUT_OBUF(m0_oper0_waddr[2]));

	IBUF QL_INST_A2F_T_4_0 (.IN_IBUF(m0_oper0_rdata[21]),.OUT_IBUF(m0_oper0_rdata_int[21]));

	IBUF QL_INST_A2F_T_4_1 (.IN_IBUF(m0_oper0_rdata[20]),.OUT_IBUF(m0_oper0_rdata_int[20]));

	IBUF QL_INST_A2F_T_4_2 (.IN_IBUF(m0_oper0_rdata[19]),.OUT_IBUF(m0_oper0_rdata_int[19]));

	IBUF QL_INST_A2F_T_4_3 (.IN_IBUF(m0_oper0_rdata[18]),.OUT_IBUF(m0_oper0_rdata_int[18]));

	IBUF QL_INST_A2F_T_4_4 (.IN_IBUF(m0_oper0_rdata[17]),.OUT_IBUF(m0_oper0_rdata_int[17]));

	IBUF QL_INST_A2F_T_4_5 (.IN_IBUF(m0_oper0_rdata[16]),.OUT_IBUF(m0_oper0_rdata_int[16]));

	IBUF QL_INST_A2F_T_4_6 (.IN_IBUF(m0_oper0_rdata[15]),.OUT_IBUF(m0_oper0_rdata_int[15]));

	IBUF QL_INST_A2F_T_4_7 (.IN_IBUF(m0_oper0_rdata[14]),.OUT_IBUF(m0_oper0_rdata_int[14]));

	OBUF QL_INST_F2A_T_5_0 (.IN_OBUF(m0_oper0_waddr_dup_0[1]),.OUT_OBUF(m0_oper0_waddr[1]));

	OBUF QL_INST_F2A_T_5_1 (.IN_OBUF(m0_oper0_waddr_dup_0[0]),.OUT_OBUF(m0_oper0_waddr[0]));

	OBUF QL_INST_F2A_T_5_2 (.IN_OBUF(m0_oper0_we_dup_0),.OUT_OBUF(m0_oper0_we));

	OBUF QL_INST_F2A_T_5_3 (.IN_OBUF(m0_oper0_raddr_dup_0[11]),.OUT_OBUF(m0_oper0_raddr[11]));

	OBUF QL_INST_F2A_T_5_4 (.IN_OBUF(m0_oper0_raddr_dup_0[10]),.OUT_OBUF(m0_oper0_raddr[10]));

	OBUF QL_INST_F2A_T_5_5 (.IN_OBUF(m0_oper0_raddr_dup_0[9]),.OUT_OBUF(m0_oper0_raddr[9]));

	OBUF QL_INST_F2A_T_5_6 (.IN_OBUF(m0_oper0_raddr_dup_0[8]),.OUT_OBUF(m0_oper0_raddr[8]));

	OBUF QL_INST_F2A_T_5_7 (.IN_OBUF(m0_oper0_raddr_dup_0[7]),.OUT_OBUF(m0_oper0_raddr[7]));

	OBUF QL_INST_F2A_T_5_8 (.IN_OBUF(m0_oper0_raddr_dup_0[6]),.OUT_OBUF(m0_oper0_raddr[6]));

	OBUF QL_INST_F2A_T_5_9 (.IN_OBUF(m0_oper0_raddr_dup_0[5]),.OUT_OBUF(m0_oper0_raddr[5]));

	OBUF QL_INST_F2A_T_5_10 (.IN_OBUF(m0_oper0_raddr_dup_0[4]),.OUT_OBUF(m0_oper0_raddr[4]));

	OBUF QL_INST_F2A_T_5_11 (.IN_OBUF(m0_oper0_raddr_dup_0[3]),.OUT_OBUF(m0_oper0_raddr[3]));

	IBUF QL_INST_A2F_T_5_0 (.IN_IBUF(m0_oper0_rdata[13]),.OUT_IBUF(m0_oper0_rdata_int[13]));

	IBUF QL_INST_A2F_T_5_1 (.IN_IBUF(m0_oper0_rdata[12]),.OUT_IBUF(m0_oper0_rdata_int[12]));

	IBUF QL_INST_A2F_T_5_2 (.IN_IBUF(m0_oper0_rdata[11]),.OUT_IBUF(m0_oper0_rdata_int[11]));

	IBUF QL_INST_A2F_T_5_3 (.IN_IBUF(m0_oper0_rdata[10]),.OUT_IBUF(m0_oper0_rdata_int[10]));

	IBUF QL_INST_A2F_T_5_4 (.IN_IBUF(m0_oper0_rdata[9]),.OUT_IBUF(m0_oper0_rdata_int[9]));

	IBUF QL_INST_A2F_T_5_5 (.IN_IBUF(m0_oper0_rdata[8]),.OUT_IBUF(m0_oper0_rdata_int[8]));

	OBUF QL_INST_F2A_T_6_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTL_6_padClk),.OUT_OBUF(m0_oper0_rclk));

	OBUF QL_INST_F2A_T_6_1 (.IN_OBUF(m0_oper0_raddr_dup_0[2]),.OUT_OBUF(m0_oper0_raddr[2]));

	OBUF QL_INST_F2A_T_6_2 (.IN_OBUF(m0_oper0_raddr_dup_0[1]),.OUT_OBUF(m0_oper0_raddr[1]));

	OBUF QL_INST_F2A_T_6_3 (.IN_OBUF(m0_oper0_raddr_dup_0[0]),.OUT_OBUF(m0_oper0_raddr[0]));

	OBUF QL_INST_F2A_T_6_4 (.IN_OBUF(m0_m0_osel_dup_0),.OUT_OBUF(m0_m0_osel));

	OBUF QL_INST_F2A_T_6_5 (.IN_OBUF(m0_m0_clken_dup_0),.OUT_OBUF(m0_m0_clken));

	OBUF QL_INST_F2A_T_6_6 (.IN_OBUF(m0_m0_outsel_dup_0[5]),.OUT_OBUF(m0_m0_outsel[5]));

	OBUF QL_INST_F2A_T_6_7 (.IN_OBUF(m0_m0_outsel_dup_0[4]),.OUT_OBUF(m0_m0_outsel[4]));

	OBUF QL_INST_F2A_T_6_8 (.IN_OBUF(m0_m0_outsel_dup_0[3]),.OUT_OBUF(m0_m0_outsel[3]));

	OBUF QL_INST_F2A_T_6_9 (.IN_OBUF(m0_m0_outsel_dup_0[2]),.OUT_OBUF(m0_m0_outsel[2]));

	OBUF QL_INST_F2A_T_6_10 (.IN_OBUF(m0_m0_outsel_dup_0[1]),.OUT_OBUF(m0_m0_outsel[1]));

	OBUF QL_INST_F2A_T_6_11 (.IN_OBUF(m0_m0_outsel_dup_0[0]),.OUT_OBUF(m0_m0_outsel[0]));

	OBUF QL_INST_F2A_T_6_12 (.IN_OBUF(m0_m0_sat_dup_0),.OUT_OBUF(m0_m0_sat));

	OBUF QL_INST_F2A_T_6_13 (.IN_OBUF(m0_m0_rnd_dup_0),.OUT_OBUF(m0_m0_rnd));

	OBUF QL_INST_F2A_T_6_14 (.IN_OBUF(m0_m0_clr_dup_0),.OUT_OBUF(m0_m0_clr));

	OBUF QL_INST_F2A_T_6_15 (.IN_OBUF(m0_oper0_rdata_int[31]),.OUT_OBUF(m0_m0_oper_in[31]));

	OBUF QL_INST_F2A_T_6_16 (.IN_OBUF(m0_oper0_rdata_int[30]),.OUT_OBUF(m0_m0_oper_in[30]));

	OBUF QL_INST_F2A_T_6_17 (.IN_OBUF(m0_oper0_rdata_int[29]),.OUT_OBUF(m0_m0_oper_in[29]));

	DBUF QL_INST_F2Adef_T_6_1 (.IN_DBUF(GND),.OUT_DBUF(m0_oper0_powerdn));

	IBUF QL_INST_A2F_T_6_0 (.IN_IBUF(m0_oper0_rdata[7]),.OUT_IBUF(m0_oper0_rdata_int[7]));

	IBUF QL_INST_A2F_T_6_1 (.IN_IBUF(m0_oper0_rdata[6]),.OUT_IBUF(m0_oper0_rdata_int[6]));

	IBUF QL_INST_A2F_T_6_2 (.IN_IBUF(m0_oper0_rdata[5]),.OUT_IBUF(m0_oper0_rdata_int[5]));

	IBUF QL_INST_A2F_T_6_3 (.IN_IBUF(m0_oper0_rdata[4]),.OUT_IBUF(m0_oper0_rdata_int[4]));

	IBUF QL_INST_A2F_T_6_4 (.IN_IBUF(m0_oper0_rdata[3]),.OUT_IBUF(m0_oper0_rdata_int[3]));

	IBUF QL_INST_A2F_T_6_5 (.IN_IBUF(m0_oper0_rdata[2]),.OUT_IBUF(m0_oper0_rdata_int[2]));

	IBUF QL_INST_A2F_T_6_6 (.IN_IBUF(m0_oper0_rdata[1]),.OUT_IBUF(m0_oper0_rdata_int[1]));

	IBUF QL_INST_A2F_T_6_7 (.IN_IBUF(m0_oper0_rdata[0]),.OUT_IBUF(m0_oper0_rdata_int[0]));

	OBUF QL_INST_F2A_T_7_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTL_7_padClk),.OUT_OBUF(m0_m0_clk));

	OBUF QL_INST_F2A_T_7_1 (.IN_OBUF(m0_oper0_rdata_int[28]),.OUT_OBUF(m0_m0_oper_in[28]));

	OBUF QL_INST_F2A_T_7_2 (.IN_OBUF(m0_oper0_rdata_int[27]),.OUT_OBUF(m0_m0_oper_in[27]));

	OBUF QL_INST_F2A_T_7_3 (.IN_OBUF(m0_oper0_rdata_int[26]),.OUT_OBUF(m0_m0_oper_in[26]));

	OBUF QL_INST_F2A_T_7_4 (.IN_OBUF(m0_oper0_rdata_int[25]),.OUT_OBUF(m0_m0_oper_in[25]));

	OBUF QL_INST_F2A_T_7_5 (.IN_OBUF(m0_oper0_rdata_int[24]),.OUT_OBUF(m0_m0_oper_in[24]));

	OBUF QL_INST_F2A_T_7_6 (.IN_OBUF(m0_oper0_rdata_int[23]),.OUT_OBUF(m0_m0_oper_in[23]));

	OBUF QL_INST_F2A_T_7_7 (.IN_OBUF(m0_oper0_rdata_int[22]),.OUT_OBUF(m0_m0_oper_in[22]));

	OBUF QL_INST_F2A_T_7_8 (.IN_OBUF(m0_oper0_rdata_int[21]),.OUT_OBUF(m0_m0_oper_in[21]));

	OBUF QL_INST_F2A_T_7_9 (.IN_OBUF(m0_oper0_rdata_int[20]),.OUT_OBUF(m0_m0_oper_in[20]));

	OBUF QL_INST_F2A_T_7_10 (.IN_OBUF(m0_oper0_rdata_int[19]),.OUT_OBUF(m0_m0_oper_in[19]));

	OBUF QL_INST_F2A_T_7_11 (.IN_OBUF(m0_oper0_rdata_int[18]),.OUT_OBUF(m0_m0_oper_in[18]));

	IBUF QL_INST_A2F_T_7_0 (.IN_IBUF(m0_m0_dataout[31]),.OUT_IBUF(m0_m0_dataout_int[31]));

	IBUF QL_INST_A2F_T_7_1 (.IN_IBUF(m0_m0_dataout[30]),.OUT_IBUF(m0_m0_dataout_int[30]));

	IBUF QL_INST_A2F_T_7_2 (.IN_IBUF(m0_m0_dataout[29]),.OUT_IBUF(m0_m0_dataout_int[29]));

	IBUF QL_INST_A2F_T_7_3 (.IN_IBUF(m0_m0_dataout[28]),.OUT_IBUF(m0_m0_dataout_int[28]));

	IBUF QL_INST_A2F_T_7_4 (.IN_IBUF(m0_m0_dataout[27]),.OUT_IBUF(m0_m0_dataout_int[27]));

	IBUF QL_INST_A2F_T_7_5 (.IN_IBUF(m0_m0_dataout[26]),.OUT_IBUF(m0_m0_dataout_int[26]));

	OBUF QL_INST_F2A_T_8_0 (.IN_OBUF(m0_oper0_rdata_int[17]),.OUT_OBUF(m0_m0_oper_in[17]));

	OBUF QL_INST_F2A_T_8_1 (.IN_OBUF(m0_oper0_rdata_int[16]),.OUT_OBUF(m0_m0_oper_in[16]));

	OBUF QL_INST_F2A_T_8_2 (.IN_OBUF(m0_oper0_rdata_int[15]),.OUT_OBUF(m0_m0_oper_in[15]));

	OBUF QL_INST_F2A_T_8_3 (.IN_OBUF(m0_oper0_rdata_int[14]),.OUT_OBUF(m0_m0_oper_in[14]));

	OBUF QL_INST_F2A_T_8_4 (.IN_OBUF(m0_oper0_rdata_int[13]),.OUT_OBUF(m0_m0_oper_in[13]));

	OBUF QL_INST_F2A_T_8_5 (.IN_OBUF(m0_oper0_rdata_int[12]),.OUT_OBUF(m0_m0_oper_in[12]));

	OBUF QL_INST_F2A_T_8_6 (.IN_OBUF(m0_oper0_rdata_int[11]),.OUT_OBUF(m0_m0_oper_in[11]));

	OBUF QL_INST_F2A_T_8_7 (.IN_OBUF(m0_oper0_rdata_int[10]),.OUT_OBUF(m0_m0_oper_in[10]));

	OBUF QL_INST_F2A_T_8_8 (.IN_OBUF(m0_oper0_rdata_int[9]),.OUT_OBUF(m0_m0_oper_in[9]));

	OBUF QL_INST_F2A_T_8_9 (.IN_OBUF(m0_oper0_rdata_int[8]),.OUT_OBUF(m0_m0_oper_in[8]));

	OBUF QL_INST_F2A_T_8_10 (.IN_OBUF(m0_oper0_rdata_int[7]),.OUT_OBUF(m0_m0_oper_in[7]));

	OBUF QL_INST_F2A_T_8_11 (.IN_OBUF(m0_oper0_rdata_int[6]),.OUT_OBUF(m0_m0_oper_in[6]));

	OBUF QL_INST_F2A_T_8_12 (.IN_OBUF(m0_oper0_rdata_int[5]),.OUT_OBUF(m0_m0_oper_in[5]));

	OBUF QL_INST_F2A_T_8_13 (.IN_OBUF(m0_oper0_rdata_int[4]),.OUT_OBUF(m0_m0_oper_in[4]));

	OBUF QL_INST_F2A_T_8_14 (.IN_OBUF(m0_oper0_rdata_int[3]),.OUT_OBUF(m0_m0_oper_in[3]));

	OBUF QL_INST_F2A_T_8_15 (.IN_OBUF(m0_oper0_rdata_int[2]),.OUT_OBUF(m0_m0_oper_in[2]));

	OBUF QL_INST_F2A_T_8_16 (.IN_OBUF(m0_oper0_rdata_int[1]),.OUT_OBUF(m0_m0_oper_in[1]));

	OBUF QL_INST_F2A_T_8_17 (.IN_OBUF(m0_oper0_rdata_int[0]),.OUT_OBUF(m0_m0_oper_in[0]));

	IBUF QL_INST_A2F_T_8_0 (.IN_IBUF(m0_m0_dataout[25]),.OUT_IBUF(m0_m0_dataout_int[25]));

	IBUF QL_INST_A2F_T_8_1 (.IN_IBUF(m0_m0_dataout[24]),.OUT_IBUF(m0_m0_dataout_int[24]));

	IBUF QL_INST_A2F_T_8_2 (.IN_IBUF(m0_m0_dataout[23]),.OUT_IBUF(m0_m0_dataout_int[23]));

	IBUF QL_INST_A2F_T_8_3 (.IN_IBUF(m0_m0_dataout[22]),.OUT_IBUF(m0_m0_dataout_int[22]));

	IBUF QL_INST_A2F_T_8_4 (.IN_IBUF(m0_m0_dataout[21]),.OUT_IBUF(m0_m0_dataout_int[21]));

	IBUF QL_INST_A2F_T_8_5 (.IN_IBUF(m0_m0_dataout[20]),.OUT_IBUF(m0_m0_dataout_int[20]));

	IBUF QL_INST_A2F_T_8_6 (.IN_IBUF(m0_m0_dataout[19]),.OUT_IBUF(m0_m0_dataout_int[19]));

	IBUF QL_INST_A2F_T_8_7 (.IN_IBUF(m0_m0_dataout[18]),.OUT_IBUF(m0_m0_dataout_int[18]));

	OBUF QL_INST_F2A_T_9_0 (.IN_OBUF(m0_m0_csel_dup_0),.OUT_OBUF(m0_m0_csel));

	OBUF QL_INST_F2A_T_9_1 (.IN_OBUF(m0_coef_rdata_int[31]),.OUT_OBUF(m0_m0_coef_in[31]));

	OBUF QL_INST_F2A_T_9_2 (.IN_OBUF(m0_coef_rdata_int[30]),.OUT_OBUF(m0_m0_coef_in[30]));

	OBUF QL_INST_F2A_T_9_3 (.IN_OBUF(m0_coef_rdata_int[29]),.OUT_OBUF(m0_m0_coef_in[29]));

	OBUF QL_INST_F2A_T_9_4 (.IN_OBUF(m0_coef_rdata_int[28]),.OUT_OBUF(m0_m0_coef_in[28]));

	OBUF QL_INST_F2A_T_9_5 (.IN_OBUF(m0_coef_rdata_int[27]),.OUT_OBUF(m0_m0_coef_in[27]));

	OBUF QL_INST_F2A_T_9_6 (.IN_OBUF(m0_coef_rdata_int[26]),.OUT_OBUF(m0_m0_coef_in[26]));

	OBUF QL_INST_F2A_T_9_7 (.IN_OBUF(m0_coef_rdata_int[25]),.OUT_OBUF(m0_m0_coef_in[25]));

	OBUF QL_INST_F2A_T_9_8 (.IN_OBUF(m0_coef_rdata_int[24]),.OUT_OBUF(m0_m0_coef_in[24]));

	OBUF QL_INST_F2A_T_9_9 (.IN_OBUF(m0_coef_rdata_int[23]),.OUT_OBUF(m0_m0_coef_in[23]));

	OBUF QL_INST_F2A_T_9_10 (.IN_OBUF(m0_coef_rdata_int[22]),.OUT_OBUF(m0_m0_coef_in[22]));

	OBUF QL_INST_F2A_T_9_11 (.IN_OBUF(m0_coef_rdata_int[21]),.OUT_OBUF(m0_m0_coef_in[21]));

	IBUF QL_INST_A2F_T_9_0 (.IN_IBUF(m0_m0_dataout[17]),.OUT_IBUF(m0_m0_dataout_int[17]));

	IBUF QL_INST_A2F_T_9_1 (.IN_IBUF(m0_m0_dataout[16]),.OUT_IBUF(m0_m0_dataout_int[16]));

	IBUF QL_INST_A2F_T_9_2 (.IN_IBUF(m0_m0_dataout[15]),.OUT_IBUF(m0_m0_dataout_int[15]));

	IBUF QL_INST_A2F_T_9_3 (.IN_IBUF(m0_m0_dataout[14]),.OUT_IBUF(m0_m0_dataout_int[14]));

	IBUF QL_INST_A2F_T_9_4 (.IN_IBUF(m0_m0_dataout[13]),.OUT_IBUF(m0_m0_dataout_int[13]));

	IBUF QL_INST_A2F_T_9_5 (.IN_IBUF(m0_m0_dataout[12]),.OUT_IBUF(m0_m0_dataout_int[12]));

	OBUF QL_INST_F2A_T_10_0 (.IN_OBUF(m0_coef_rdata_int[20]),.OUT_OBUF(m0_m0_coef_in[20]));

	OBUF QL_INST_F2A_T_10_1 (.IN_OBUF(m0_coef_rdata_int[19]),.OUT_OBUF(m0_m0_coef_in[19]));

	OBUF QL_INST_F2A_T_10_2 (.IN_OBUF(m0_coef_rdata_int[18]),.OUT_OBUF(m0_m0_coef_in[18]));

	OBUF QL_INST_F2A_T_10_3 (.IN_OBUF(m0_coef_rdata_int[17]),.OUT_OBUF(m0_m0_coef_in[17]));

	OBUF QL_INST_F2A_T_10_4 (.IN_OBUF(m0_coef_rdata_int[16]),.OUT_OBUF(m0_m0_coef_in[16]));

	OBUF QL_INST_F2A_T_10_5 (.IN_OBUF(m0_coef_rdata_int[15]),.OUT_OBUF(m0_m0_coef_in[15]));

	OBUF QL_INST_F2A_T_10_6 (.IN_OBUF(m0_coef_rdata_int[14]),.OUT_OBUF(m0_m0_coef_in[14]));

	OBUF QL_INST_F2A_T_10_7 (.IN_OBUF(m0_coef_rdata_int[13]),.OUT_OBUF(m0_m0_coef_in[13]));

	OBUF QL_INST_F2A_T_10_8 (.IN_OBUF(m0_coef_rdata_int[12]),.OUT_OBUF(m0_m0_coef_in[12]));

	OBUF QL_INST_F2A_T_10_9 (.IN_OBUF(m0_coef_rdata_int[11]),.OUT_OBUF(m0_m0_coef_in[11]));

	OBUF QL_INST_F2A_T_10_10 (.IN_OBUF(m0_coef_rdata_int[10]),.OUT_OBUF(m0_m0_coef_in[10]));

	OBUF QL_INST_F2A_T_10_11 (.IN_OBUF(m0_coef_rdata_int[9]),.OUT_OBUF(m0_m0_coef_in[9]));

	OBUF QL_INST_F2A_T_10_12 (.IN_OBUF(m0_coef_rdata_int[8]),.OUT_OBUF(m0_m0_coef_in[8]));

	OBUF QL_INST_F2A_T_10_13 (.IN_OBUF(m0_coef_rdata_int[7]),.OUT_OBUF(m0_m0_coef_in[7]));

	OBUF QL_INST_F2A_T_10_14 (.IN_OBUF(m0_coef_rdata_int[6]),.OUT_OBUF(m0_m0_coef_in[6]));

	OBUF QL_INST_F2A_T_10_15 (.IN_OBUF(m0_coef_rdata_int[5]),.OUT_OBUF(m0_m0_coef_in[5]));

	OBUF QL_INST_F2A_T_10_16 (.IN_OBUF(m0_coef_rdata_int[4]),.OUT_OBUF(m0_m0_coef_in[4]));

	OBUF QL_INST_F2A_T_10_17 (.IN_OBUF(m0_coef_rdata_int[3]),.OUT_OBUF(m0_m0_coef_in[3]));

	IBUF QL_INST_A2F_T_10_0 (.IN_IBUF(m0_m0_dataout[11]),.OUT_IBUF(m0_m0_dataout_int[11]));

	IBUF QL_INST_A2F_T_10_1 (.IN_IBUF(m0_m0_dataout[10]),.OUT_IBUF(m0_m0_dataout_int[10]));

	IBUF QL_INST_A2F_T_10_2 (.IN_IBUF(m0_m0_dataout[9]),.OUT_IBUF(m0_m0_dataout_int[9]));

	IBUF QL_INST_A2F_T_10_3 (.IN_IBUF(m0_m0_dataout[8]),.OUT_IBUF(m0_m0_dataout_int[8]));

	IBUF QL_INST_A2F_T_10_4 (.IN_IBUF(m0_m0_dataout[7]),.OUT_IBUF(m0_m0_dataout_int[7]));

	IBUF QL_INST_A2F_T_10_5 (.IN_IBUF(m0_m0_dataout[6]),.OUT_IBUF(m0_m0_dataout_int[6]));

	IBUF QL_INST_A2F_T_10_6 (.IN_IBUF(m0_m0_dataout[5]),.OUT_IBUF(m0_m0_dataout_int[5]));

	IBUF QL_INST_A2F_T_10_7 (.IN_IBUF(m0_m0_dataout[4]),.OUT_IBUF(m0_m0_dataout_int[4]));

	OBUF QL_INST_F2A_T_11_0 (.IN_OBUF(m0_coef_rdata_int[2]),.OUT_OBUF(m0_m0_coef_in[2]));

	OBUF QL_INST_F2A_T_11_1 (.IN_OBUF(m0_coef_rdata_int[1]),.OUT_OBUF(m0_m0_coef_in[1]));

	OBUF QL_INST_F2A_T_11_2 (.IN_OBUF(m0_coef_rdata_int[0]),.OUT_OBUF(m0_m0_coef_in[0]));

	OBUF QL_INST_F2A_T_11_3 (.IN_OBUF(m0_m0_mode_dup_0[1]),.OUT_OBUF(m0_m0_mode[1]));

	OBUF QL_INST_F2A_T_11_4 (.IN_OBUF(m0_m0_mode_dup_0[0]),.OUT_OBUF(m0_m0_mode[0]));

	OBUF QL_INST_F2A_T_11_5 (.IN_OBUF(m0_m0_tc_dup_0),.OUT_OBUF(m0_m0_tc));

	OBUF QL_INST_F2A_T_11_6 (.IN_OBUF(m0_m0_reset_dup_0),.OUT_OBUF(m0_m0_reset));

	OBUF QL_INST_F2A_T_11_7 (.IN_OBUF(m0_coef_wdata_dup_0[31]),.OUT_OBUF(m0_coef_wdata[31]));

	OBUF QL_INST_F2A_T_11_8 (.IN_OBUF(m0_coef_wdata_dup_0[30]),.OUT_OBUF(m0_coef_wdata[30]));

	OBUF QL_INST_F2A_T_11_9 (.IN_OBUF(m0_coef_wdata_dup_0[29]),.OUT_OBUF(m0_coef_wdata[29]));

	OBUF QL_INST_F2A_T_11_10 (.IN_OBUF(m0_coef_wdata_dup_0[28]),.OUT_OBUF(m0_coef_wdata[28]));

	OBUF QL_INST_F2A_T_11_11 (.IN_OBUF(m0_coef_wdata_dup_0[27]),.OUT_OBUF(m0_coef_wdata[27]));

	IBUF QL_INST_A2F_T_11_0 (.IN_IBUF(m0_m0_dataout[3]),.OUT_IBUF(m0_m0_dataout_int[3]));

	IBUF QL_INST_A2F_T_11_1 (.IN_IBUF(m0_m0_dataout[2]),.OUT_IBUF(m0_m0_dataout_int[2]));

	IBUF QL_INST_A2F_T_11_2 (.IN_IBUF(m0_m0_dataout[1]),.OUT_IBUF(m0_m0_dataout_int[1]));

	IBUF QL_INST_A2F_T_11_3 (.IN_IBUF(m0_m0_dataout[0]),.OUT_IBUF(m0_m0_dataout_int[0]));

	IBUF QL_INST_A2F_T_11_4 (.IN_IBUF(m0_coef_rdata[31]),.OUT_IBUF(m0_coef_rdata_int[31]));

	IBUF QL_INST_A2F_T_11_5 (.IN_IBUF(m0_coef_rdata[30]),.OUT_IBUF(m0_coef_rdata_int[30]));

	OBUF QL_INST_F2A_T_12_0 (.IN_OBUF(m0_coef_wdata_dup_0[26]),.OUT_OBUF(m0_coef_wdata[26]));

	OBUF QL_INST_F2A_T_12_1 (.IN_OBUF(m0_coef_wdata_dup_0[25]),.OUT_OBUF(m0_coef_wdata[25]));

	OBUF QL_INST_F2A_T_12_2 (.IN_OBUF(m0_coef_wdata_dup_0[24]),.OUT_OBUF(m0_coef_wdata[24]));

	OBUF QL_INST_F2A_T_12_3 (.IN_OBUF(m0_coef_wdata_dup_0[23]),.OUT_OBUF(m0_coef_wdata[23]));

	OBUF QL_INST_F2A_T_12_4 (.IN_OBUF(m0_coef_wdata_dup_0[22]),.OUT_OBUF(m0_coef_wdata[22]));

	OBUF QL_INST_F2A_T_12_5 (.IN_OBUF(m0_coef_wdata_dup_0[21]),.OUT_OBUF(m0_coef_wdata[21]));

	OBUF QL_INST_F2A_T_12_6 (.IN_OBUF(m0_coef_wdata_dup_0[20]),.OUT_OBUF(m0_coef_wdata[20]));

	OBUF QL_INST_F2A_T_12_7 (.IN_OBUF(m0_coef_wdata_dup_0[19]),.OUT_OBUF(m0_coef_wdata[19]));

	OBUF QL_INST_F2A_T_12_8 (.IN_OBUF(m0_coef_wdata_dup_0[18]),.OUT_OBUF(m0_coef_wdata[18]));

	OBUF QL_INST_F2A_T_12_9 (.IN_OBUF(m0_coef_wdata_dup_0[17]),.OUT_OBUF(m0_coef_wdata[17]));

	OBUF QL_INST_F2A_T_12_10 (.IN_OBUF(m0_coef_wdata_dup_0[16]),.OUT_OBUF(m0_coef_wdata[16]));

	OBUF QL_INST_F2A_T_12_11 (.IN_OBUF(m0_coef_wdata_dup_0[15]),.OUT_OBUF(m0_coef_wdata[15]));

	OBUF QL_INST_F2A_T_12_12 (.IN_OBUF(m0_coef_wdata_dup_0[14]),.OUT_OBUF(m0_coef_wdata[14]));

	OBUF QL_INST_F2A_T_12_13 (.IN_OBUF(m0_coef_wdata_dup_0[13]),.OUT_OBUF(m0_coef_wdata[13]));

	OBUF QL_INST_F2A_T_12_14 (.IN_OBUF(m0_coef_wdata_dup_0[12]),.OUT_OBUF(m0_coef_wdata[12]));

	OBUF QL_INST_F2A_T_12_15 (.IN_OBUF(m0_coef_wdata_dup_0[11]),.OUT_OBUF(m0_coef_wdata[11]));

	OBUF QL_INST_F2A_T_12_16 (.IN_OBUF(m0_coef_wdata_dup_0[10]),.OUT_OBUF(m0_coef_wdata[10]));

	OBUF QL_INST_F2A_T_12_17 (.IN_OBUF(m0_coef_wdata_dup_0[9]),.OUT_OBUF(m0_coef_wdata[9]));

	IBUF QL_INST_A2F_T_12_0 (.IN_IBUF(m0_coef_rdata[29]),.OUT_IBUF(m0_coef_rdata_int[29]));

	IBUF QL_INST_A2F_T_12_1 (.IN_IBUF(m0_coef_rdata[28]),.OUT_IBUF(m0_coef_rdata_int[28]));

	IBUF QL_INST_A2F_T_12_2 (.IN_IBUF(m0_coef_rdata[27]),.OUT_IBUF(m0_coef_rdata_int[27]));

	IBUF QL_INST_A2F_T_12_3 (.IN_IBUF(m0_coef_rdata[26]),.OUT_IBUF(m0_coef_rdata_int[26]));

	IBUF QL_INST_A2F_T_12_4 (.IN_IBUF(m0_coef_rdata[25]),.OUT_IBUF(m0_coef_rdata_int[25]));

	IBUF QL_INST_A2F_T_12_5 (.IN_IBUF(m0_coef_rdata[24]),.OUT_IBUF(m0_coef_rdata_int[24]));

	IBUF QL_INST_A2F_T_12_6 (.IN_IBUF(m0_coef_rdata[23]),.OUT_IBUF(m0_coef_rdata_int[23]));

	IBUF QL_INST_A2F_T_12_7 (.IN_IBUF(m0_coef_rdata[22]),.OUT_IBUF(m0_coef_rdata_int[22]));

	OBUF QL_INST_F2A_T_13_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTR_13_padClk),.OUT_OBUF(m0_coef_wclk));

	OBUF QL_INST_F2A_T_13_1 (.IN_OBUF(m0_coef_wdata_dup_0[8]),.OUT_OBUF(m0_coef_wdata[8]));

	OBUF QL_INST_F2A_T_13_2 (.IN_OBUF(m0_coef_wdata_dup_0[7]),.OUT_OBUF(m0_coef_wdata[7]));

	OBUF QL_INST_F2A_T_13_3 (.IN_OBUF(m0_coef_wdata_dup_0[6]),.OUT_OBUF(m0_coef_wdata[6]));

	OBUF QL_INST_F2A_T_13_4 (.IN_OBUF(m0_coef_wdata_dup_0[5]),.OUT_OBUF(m0_coef_wdata[5]));

	OBUF QL_INST_F2A_T_13_5 (.IN_OBUF(m0_coef_wdata_dup_0[4]),.OUT_OBUF(m0_coef_wdata[4]));

	OBUF QL_INST_F2A_T_13_6 (.IN_OBUF(m0_coef_wdata_dup_0[3]),.OUT_OBUF(m0_coef_wdata[3]));

	OBUF QL_INST_F2A_T_13_7 (.IN_OBUF(m0_coef_wdata_dup_0[2]),.OUT_OBUF(m0_coef_wdata[2]));

	OBUF QL_INST_F2A_T_13_8 (.IN_OBUF(m0_coef_wdata_dup_0[1]),.OUT_OBUF(m0_coef_wdata[1]));

	OBUF QL_INST_F2A_T_13_9 (.IN_OBUF(m0_coef_wdata_dup_0[0]),.OUT_OBUF(m0_coef_wdata[0]));

	OBUF QL_INST_F2A_T_13_10 (.IN_OBUF(m0_coef_waddr_dup_0[11]),.OUT_OBUF(m0_coef_waddr[11]));

	OBUF QL_INST_F2A_T_13_11 (.IN_OBUF(m0_coef_waddr_dup_0[10]),.OUT_OBUF(m0_coef_waddr[10]));

	DBUF QL_INST_F2Adef_T_13_0 (.IN_DBUF(GND),.OUT_DBUF(m0_coef_powerdn));

	IBUF QL_INST_A2F_T_13_0 (.IN_IBUF(m0_coef_rdata[21]),.OUT_IBUF(m0_coef_rdata_int[21]));

	IBUF QL_INST_A2F_T_13_1 (.IN_IBUF(m0_coef_rdata[20]),.OUT_IBUF(m0_coef_rdata_int[20]));

	IBUF QL_INST_A2F_T_13_2 (.IN_IBUF(m0_coef_rdata[19]),.OUT_IBUF(m0_coef_rdata_int[19]));

	IBUF QL_INST_A2F_T_13_3 (.IN_IBUF(m0_coef_rdata[18]),.OUT_IBUF(m0_coef_rdata_int[18]));

	IBUF QL_INST_A2F_T_13_4 (.IN_IBUF(m0_coef_rdata[17]),.OUT_IBUF(m0_coef_rdata_int[17]));

	IBUF QL_INST_A2F_T_13_5 (.IN_IBUF(m0_coef_rdata[16]),.OUT_IBUF(m0_coef_rdata_int[16]));

	OBUF QL_INST_F2A_T_14_0 (.IN_OBUF(m0_coef_waddr_dup_0[9]),.OUT_OBUF(m0_coef_waddr[9]));

	OBUF QL_INST_F2A_T_14_1 (.IN_OBUF(m0_coef_waddr_dup_0[8]),.OUT_OBUF(m0_coef_waddr[8]));

	OBUF QL_INST_F2A_T_14_2 (.IN_OBUF(m0_coef_waddr_dup_0[7]),.OUT_OBUF(m0_coef_waddr[7]));

	OBUF QL_INST_F2A_T_14_3 (.IN_OBUF(m0_coef_waddr_dup_0[6]),.OUT_OBUF(m0_coef_waddr[6]));

	OBUF QL_INST_F2A_T_14_4 (.IN_OBUF(m0_coef_waddr_dup_0[5]),.OUT_OBUF(m0_coef_waddr[5]));

	OBUF QL_INST_F2A_T_14_5 (.IN_OBUF(m0_coef_waddr_dup_0[4]),.OUT_OBUF(m0_coef_waddr[4]));

	OBUF QL_INST_F2A_T_14_6 (.IN_OBUF(m0_coef_waddr_dup_0[3]),.OUT_OBUF(m0_coef_waddr[3]));

	OBUF QL_INST_F2A_T_14_7 (.IN_OBUF(m0_coef_waddr_dup_0[2]),.OUT_OBUF(m0_coef_waddr[2]));

	OBUF QL_INST_F2A_T_14_8 (.IN_OBUF(m0_coef_waddr_dup_0[1]),.OUT_OBUF(m0_coef_waddr[1]));

	OBUF QL_INST_F2A_T_14_9 (.IN_OBUF(m0_coef_waddr_dup_0[0]),.OUT_OBUF(m0_coef_waddr[0]));

	OBUF QL_INST_F2A_T_14_10 (.IN_OBUF(m0_coef_we_dup_0),.OUT_OBUF(m0_coef_we));

	OBUF QL_INST_F2A_T_14_11 (.IN_OBUF(m0_coef_wdsel_dup_0),.OUT_OBUF(m0_coef_wdsel));

	OBUF QL_INST_F2A_T_14_12 (.IN_OBUF(m0_coef_rmode_dup_0[1]),.OUT_OBUF(m0_coef_rmode[1]));

	OBUF QL_INST_F2A_T_14_13 (.IN_OBUF(m0_coef_rmode_dup_0[0]),.OUT_OBUF(m0_coef_rmode[0]));

	OBUF QL_INST_F2A_T_14_14 (.IN_OBUF(m0_coef_raddr_dup_0[11]),.OUT_OBUF(m0_coef_raddr[11]));

	OBUF QL_INST_F2A_T_14_15 (.IN_OBUF(m0_coef_raddr_dup_0[10]),.OUT_OBUF(m0_coef_raddr[10]));

	OBUF QL_INST_F2A_T_14_16 (.IN_OBUF(m0_coef_raddr_dup_0[9]),.OUT_OBUF(m0_coef_raddr[9]));

	OBUF QL_INST_F2A_T_14_17 (.IN_OBUF(m0_coef_raddr_dup_0[8]),.OUT_OBUF(m0_coef_raddr[8]));

	IBUF QL_INST_A2F_T_14_0 (.IN_IBUF(m0_coef_rdata[15]),.OUT_IBUF(m0_coef_rdata_int[15]));

	IBUF QL_INST_A2F_T_14_1 (.IN_IBUF(m0_coef_rdata[14]),.OUT_IBUF(m0_coef_rdata_int[14]));

	IBUF QL_INST_A2F_T_14_2 (.IN_IBUF(m0_coef_rdata[13]),.OUT_IBUF(m0_coef_rdata_int[13]));

	IBUF QL_INST_A2F_T_14_3 (.IN_IBUF(m0_coef_rdata[12]),.OUT_IBUF(m0_coef_rdata_int[12]));

	IBUF QL_INST_A2F_T_14_4 (.IN_IBUF(m0_coef_rdata[11]),.OUT_IBUF(m0_coef_rdata_int[11]));

	IBUF QL_INST_A2F_T_14_5 (.IN_IBUF(m0_coef_rdata[10]),.OUT_IBUF(m0_coef_rdata_int[10]));

	IBUF QL_INST_A2F_T_14_6 (.IN_IBUF(m0_coef_rdata[9]),.OUT_IBUF(m0_coef_rdata_int[9]));

	IBUF QL_INST_A2F_T_14_7 (.IN_IBUF(m0_coef_rdata[8]),.OUT_IBUF(m0_coef_rdata_int[8]));

	OBUF QL_INST_F2A_T_15_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTR_15_padClk),.OUT_OBUF(m0_coef_rclk));

	OBUF QL_INST_F2A_T_15_1 (.IN_OBUF(m0_coef_raddr_dup_0[7]),.OUT_OBUF(m0_coef_raddr[7]));

	OBUF QL_INST_F2A_T_15_2 (.IN_OBUF(m0_coef_raddr_dup_0[6]),.OUT_OBUF(m0_coef_raddr[6]));

	OBUF QL_INST_F2A_T_15_3 (.IN_OBUF(m0_coef_raddr_dup_0[5]),.OUT_OBUF(m0_coef_raddr[5]));

	OBUF QL_INST_F2A_T_15_4 (.IN_OBUF(m0_coef_raddr_dup_0[4]),.OUT_OBUF(m0_coef_raddr[4]));

	OBUF QL_INST_F2A_T_15_5 (.IN_OBUF(m0_coef_raddr_dup_0[3]),.OUT_OBUF(m0_coef_raddr[3]));

	OBUF QL_INST_F2A_T_15_6 (.IN_OBUF(m0_coef_raddr_dup_0[2]),.OUT_OBUF(m0_coef_raddr[2]));

	OBUF QL_INST_F2A_T_15_7 (.IN_OBUF(m0_coef_raddr_dup_0[1]),.OUT_OBUF(m0_coef_raddr[1]));

	OBUF QL_INST_F2A_T_15_8 (.IN_OBUF(m0_coef_raddr_dup_0[0]),.OUT_OBUF(m0_coef_raddr[0]));

	OBUF QL_INST_F2A_T_15_9 (.IN_OBUF(m0_coef_wmode_dup_0[1]),.OUT_OBUF(m0_coef_wmode[1]));

	OBUF QL_INST_F2A_T_15_10 (.IN_OBUF(m0_coef_wmode_dup_0[0]),.OUT_OBUF(m0_coef_wmode[0]));

	IBUF QL_INST_A2F_T_15_0 (.IN_IBUF(m0_coef_rdata[7]),.OUT_IBUF(m0_coef_rdata_int[7]));

	IBUF QL_INST_A2F_T_15_1 (.IN_IBUF(m0_coef_rdata[6]),.OUT_IBUF(m0_coef_rdata_int[6]));

	IBUF QL_INST_A2F_T_15_2 (.IN_IBUF(m0_coef_rdata[5]),.OUT_IBUF(m0_coef_rdata_int[5]));

	IBUF QL_INST_A2F_T_15_3 (.IN_IBUF(m0_coef_rdata[4]),.OUT_IBUF(m0_coef_rdata_int[4]));

	IBUF QL_INST_A2F_T_15_4 (.IN_IBUF(m0_coef_rdata[3]),.OUT_IBUF(m0_coef_rdata_int[3]));

	IBUF QL_INST_A2F_T_15_5 (.IN_IBUF(m0_coef_rdata[2]),.OUT_IBUF(m0_coef_rdata_int[2]));

	IBUF QL_INST_A2F_T_16_0 (.IN_IBUF(m0_coef_rdata[1]),.OUT_IBUF(m0_coef_rdata_int[1]));

	IBUF QL_INST_A2F_T_16_1 (.IN_IBUF(m0_coef_rdata[0]),.OUT_IBUF(m0_coef_rdata_int[0]));

	OBUF QL_INST_F2A_T_18_8 (.IN_OBUF(m0_m1_outsel_dup_0[5]),.OUT_OBUF(m0_m1_outsel[5]));

	OBUF QL_INST_F2A_T_18_9 (.IN_OBUF(m0_m1_outsel_dup_0[4]),.OUT_OBUF(m0_m1_outsel[4]));

	OBUF QL_INST_F2A_T_18_10 (.IN_OBUF(m0_m1_outsel_dup_0[3]),.OUT_OBUF(m0_m1_outsel[3]));

	OBUF QL_INST_F2A_T_18_11 (.IN_OBUF(m0_m1_outsel_dup_0[2]),.OUT_OBUF(m0_m1_outsel[2]));

	OBUF QL_INST_F2A_T_18_12 (.IN_OBUF(m0_m1_outsel_dup_0[1]),.OUT_OBUF(m0_m1_outsel[1]));

	OBUF QL_INST_F2A_T_18_13 (.IN_OBUF(m0_m1_outsel_dup_0[0]),.OUT_OBUF(m0_m1_outsel[0]));

	OBUF QL_INST_F2A_T_18_14 (.IN_OBUF(m0_m1_sat_dup_0),.OUT_OBUF(m0_m1_sat));

	OBUF QL_INST_F2A_T_18_15 (.IN_OBUF(m0_m1_rnd_dup_0),.OUT_OBUF(m0_m1_rnd));

	OBUF QL_INST_F2A_T_18_16 (.IN_OBUF(m0_m1_clr_dup_0),.OUT_OBUF(m0_m1_clr));

	OBUF QL_INST_F2A_T_18_17 (.IN_OBUF(m0_m1_clken_dup_0),.OUT_OBUF(m0_m1_clken));

	IBUF QL_INST_A2F_T_18_0 (.IN_IBUF(m0_m1_dataout[31]),.OUT_IBUF(m0_m1_dataout_int[31]));

	IBUF QL_INST_A2F_T_18_1 (.IN_IBUF(m0_m1_dataout[30]),.OUT_IBUF(m0_m1_dataout_int[30]));

	IBUF QL_INST_A2F_T_18_2 (.IN_IBUF(m0_m1_dataout[29]),.OUT_IBUF(m0_m1_dataout_int[29]));

	IBUF QL_INST_A2F_T_18_3 (.IN_IBUF(m0_m1_dataout[28]),.OUT_IBUF(m0_m1_dataout_int[28]));

	IBUF QL_INST_A2F_T_18_4 (.IN_IBUF(m0_m1_dataout[27]),.OUT_IBUF(m0_m1_dataout_int[27]));

	IBUF QL_INST_A2F_T_18_5 (.IN_IBUF(m0_m1_dataout[26]),.OUT_IBUF(m0_m1_dataout_int[26]));

	IBUF QL_INST_A2F_T_18_6 (.IN_IBUF(m0_m1_dataout[25]),.OUT_IBUF(m0_m1_dataout_int[25]));

	IBUF QL_INST_A2F_T_18_7 (.IN_IBUF(m0_m1_dataout[24]),.OUT_IBUF(m0_m1_dataout_int[24]));

	OBUF QL_INST_F2A_T_19_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTL_19_padClk),.OUT_OBUF(m0_m1_clk));

	OBUF QL_INST_F2A_T_19_1 (.IN_OBUF(m0_m1_osel_dup_0),.OUT_OBUF(m0_m1_osel));

	OBUF QL_INST_F2A_T_19_2 (.IN_OBUF(m0_m1_tc_dup_0),.OUT_OBUF(m0_m1_tc));

	OBUF QL_INST_F2A_T_19_3 (.IN_OBUF(m0_m1_reset_dup_0),.OUT_OBUF(m0_m1_reset));

	OBUF QL_INST_F2A_T_19_4 (.IN_OBUF(m0_coef_rdata_int[31]),.OUT_OBUF(m0_m1_coef_in[31]));

	OBUF QL_INST_F2A_T_19_5 (.IN_OBUF(m0_coef_rdata_int[30]),.OUT_OBUF(m0_m1_coef_in[30]));

	OBUF QL_INST_F2A_T_19_6 (.IN_OBUF(m0_coef_rdata_int[29]),.OUT_OBUF(m0_m1_coef_in[29]));

	OBUF QL_INST_F2A_T_19_7 (.IN_OBUF(m0_coef_rdata_int[28]),.OUT_OBUF(m0_m1_coef_in[28]));

	OBUF QL_INST_F2A_T_19_8 (.IN_OBUF(m0_coef_rdata_int[27]),.OUT_OBUF(m0_m1_coef_in[27]));

	OBUF QL_INST_F2A_T_19_9 (.IN_OBUF(m0_coef_rdata_int[26]),.OUT_OBUF(m0_m1_coef_in[26]));

	OBUF QL_INST_F2A_T_19_10 (.IN_OBUF(m0_coef_rdata_int[25]),.OUT_OBUF(m0_m1_coef_in[25]));

	OBUF QL_INST_F2A_T_19_11 (.IN_OBUF(m0_coef_rdata_int[24]),.OUT_OBUF(m0_m1_coef_in[24]));

	IBUF QL_INST_A2F_T_19_0 (.IN_IBUF(m0_m1_dataout[23]),.OUT_IBUF(m0_m1_dataout_int[23]));

	IBUF QL_INST_A2F_T_19_1 (.IN_IBUF(m0_m1_dataout[22]),.OUT_IBUF(m0_m1_dataout_int[22]));

	IBUF QL_INST_A2F_T_19_2 (.IN_IBUF(m0_m1_dataout[21]),.OUT_IBUF(m0_m1_dataout_int[21]));

	IBUF QL_INST_A2F_T_19_3 (.IN_IBUF(m0_m1_dataout[20]),.OUT_IBUF(m0_m1_dataout_int[20]));

	IBUF QL_INST_A2F_T_19_4 (.IN_IBUF(m0_m1_dataout[19]),.OUT_IBUF(m0_m1_dataout_int[19]));

	IBUF QL_INST_A2F_T_19_5 (.IN_IBUF(m0_m1_dataout[18]),.OUT_IBUF(m0_m1_dataout_int[18]));

	OBUF QL_INST_F2A_T_20_0 (.IN_OBUF(m0_coef_rdata_int[23]),.OUT_OBUF(m0_m1_coef_in[23]));

	OBUF QL_INST_F2A_T_20_1 (.IN_OBUF(m0_coef_rdata_int[22]),.OUT_OBUF(m0_m1_coef_in[22]));

	OBUF QL_INST_F2A_T_20_2 (.IN_OBUF(m0_coef_rdata_int[21]),.OUT_OBUF(m0_m1_coef_in[21]));

	OBUF QL_INST_F2A_T_20_3 (.IN_OBUF(m0_coef_rdata_int[20]),.OUT_OBUF(m0_m1_coef_in[20]));

	OBUF QL_INST_F2A_T_20_4 (.IN_OBUF(m0_coef_rdata_int[19]),.OUT_OBUF(m0_m1_coef_in[19]));

	OBUF QL_INST_F2A_T_20_5 (.IN_OBUF(m0_coef_rdata_int[18]),.OUT_OBUF(m0_m1_coef_in[18]));

	OBUF QL_INST_F2A_T_20_6 (.IN_OBUF(m0_coef_rdata_int[17]),.OUT_OBUF(m0_m1_coef_in[17]));

	OBUF QL_INST_F2A_T_20_7 (.IN_OBUF(m0_coef_rdata_int[16]),.OUT_OBUF(m0_m1_coef_in[16]));

	OBUF QL_INST_F2A_T_20_8 (.IN_OBUF(m0_coef_rdata_int[15]),.OUT_OBUF(m0_m1_coef_in[15]));

	OBUF QL_INST_F2A_T_20_9 (.IN_OBUF(m0_coef_rdata_int[14]),.OUT_OBUF(m0_m1_coef_in[14]));

	OBUF QL_INST_F2A_T_20_10 (.IN_OBUF(m0_coef_rdata_int[13]),.OUT_OBUF(m0_m1_coef_in[13]));

	OBUF QL_INST_F2A_T_20_11 (.IN_OBUF(m0_coef_rdata_int[12]),.OUT_OBUF(m0_m1_coef_in[12]));

	OBUF QL_INST_F2A_T_20_12 (.IN_OBUF(m0_coef_rdata_int[11]),.OUT_OBUF(m0_m1_coef_in[11]));

	OBUF QL_INST_F2A_T_20_13 (.IN_OBUF(m0_coef_rdata_int[10]),.OUT_OBUF(m0_m1_coef_in[10]));

	OBUF QL_INST_F2A_T_20_14 (.IN_OBUF(m0_coef_rdata_int[9]),.OUT_OBUF(m0_m1_coef_in[9]));

	OBUF QL_INST_F2A_T_20_15 (.IN_OBUF(m0_coef_rdata_int[8]),.OUT_OBUF(m0_m1_coef_in[8]));

	OBUF QL_INST_F2A_T_20_16 (.IN_OBUF(m0_coef_rdata_int[7]),.OUT_OBUF(m0_m1_coef_in[7]));

	OBUF QL_INST_F2A_T_20_17 (.IN_OBUF(m0_coef_rdata_int[6]),.OUT_OBUF(m0_m1_coef_in[6]));

	IBUF QL_INST_A2F_T_20_0 (.IN_IBUF(m0_m1_dataout[17]),.OUT_IBUF(m0_m1_dataout_int[17]));

	IBUF QL_INST_A2F_T_20_1 (.IN_IBUF(m0_m1_dataout[16]),.OUT_IBUF(m0_m1_dataout_int[16]));

	IBUF QL_INST_A2F_T_20_2 (.IN_IBUF(m0_m1_dataout[15]),.OUT_IBUF(m0_m1_dataout_int[15]));

	IBUF QL_INST_A2F_T_20_3 (.IN_IBUF(m0_m1_dataout[14]),.OUT_IBUF(m0_m1_dataout_int[14]));

	IBUF QL_INST_A2F_T_20_4 (.IN_IBUF(m0_m1_dataout[13]),.OUT_IBUF(m0_m1_dataout_int[13]));

	IBUF QL_INST_A2F_T_20_5 (.IN_IBUF(m0_m1_dataout[12]),.OUT_IBUF(m0_m1_dataout_int[12]));

	IBUF QL_INST_A2F_T_20_6 (.IN_IBUF(m0_m1_dataout[11]),.OUT_IBUF(m0_m1_dataout_int[11]));

	OBUF QL_INST_F2A_T_21_0 (.IN_OBUF(m0_coef_rdata_int[5]),.OUT_OBUF(m0_m1_coef_in[5]));

	OBUF QL_INST_F2A_T_21_1 (.IN_OBUF(m0_coef_rdata_int[4]),.OUT_OBUF(m0_m1_coef_in[4]));

	OBUF QL_INST_F2A_T_21_2 (.IN_OBUF(m0_coef_rdata_int[3]),.OUT_OBUF(m0_m1_coef_in[3]));

	OBUF QL_INST_F2A_T_21_3 (.IN_OBUF(m0_coef_rdata_int[2]),.OUT_OBUF(m0_m1_coef_in[2]));

	OBUF QL_INST_F2A_T_21_4 (.IN_OBUF(m0_coef_rdata_int[1]),.OUT_OBUF(m0_m1_coef_in[1]));

	OBUF QL_INST_F2A_T_21_5 (.IN_OBUF(m0_coef_rdata_int[0]),.OUT_OBUF(m0_m1_coef_in[0]));

	OBUF QL_INST_F2A_T_21_6 (.IN_OBUF(m0_m1_mode_dup_0[1]),.OUT_OBUF(m0_m1_mode[1]));

	OBUF QL_INST_F2A_T_21_7 (.IN_OBUF(m0_m1_csel_dup_0),.OUT_OBUF(m0_m1_csel));

	OBUF QL_INST_F2A_T_21_8 (.IN_OBUF(m0_m1_mode_dup_0[0]),.OUT_OBUF(m0_m1_mode[0]));

	OBUF QL_INST_F2A_T_21_9 (.IN_OBUF(m0_oper1_rdata_int[31]),.OUT_OBUF(m0_m1_oper_in[31]));

	OBUF QL_INST_F2A_T_21_10 (.IN_OBUF(m0_oper1_rdata_int[30]),.OUT_OBUF(m0_m1_oper_in[30]));

	OBUF QL_INST_F2A_T_21_11 (.IN_OBUF(m0_oper1_rdata_int[29]),.OUT_OBUF(m0_m1_oper_in[29]));

	IBUF QL_INST_A2F_T_21_0 (.IN_IBUF(m0_m1_dataout[10]),.OUT_IBUF(m0_m1_dataout_int[10]));

	IBUF QL_INST_A2F_T_21_1 (.IN_IBUF(m0_m1_dataout[9]),.OUT_IBUF(m0_m1_dataout_int[9]));

	IBUF QL_INST_A2F_T_21_2 (.IN_IBUF(m0_m1_dataout[8]),.OUT_IBUF(m0_m1_dataout_int[8]));

	IBUF QL_INST_A2F_T_21_3 (.IN_IBUF(m0_m1_dataout[7]),.OUT_IBUF(m0_m1_dataout_int[7]));

	IBUF QL_INST_A2F_T_21_4 (.IN_IBUF(m0_m1_dataout[6]),.OUT_IBUF(m0_m1_dataout_int[6]));

	IBUF QL_INST_A2F_T_21_5 (.IN_IBUF(m0_m1_dataout[5]),.OUT_IBUF(m0_m1_dataout_int[5]));

	OBUF QL_INST_F2A_T_22_0 (.IN_OBUF(m0_oper1_rdata_int[28]),.OUT_OBUF(m0_m1_oper_in[28]));

	OBUF QL_INST_F2A_T_22_1 (.IN_OBUF(m0_oper1_rdata_int[27]),.OUT_OBUF(m0_m1_oper_in[27]));

	OBUF QL_INST_F2A_T_22_2 (.IN_OBUF(m0_oper1_rdata_int[26]),.OUT_OBUF(m0_m1_oper_in[26]));

	OBUF QL_INST_F2A_T_22_3 (.IN_OBUF(m0_oper1_rdata_int[25]),.OUT_OBUF(m0_m1_oper_in[25]));

	OBUF QL_INST_F2A_T_22_4 (.IN_OBUF(m0_oper1_rdata_int[24]),.OUT_OBUF(m0_m1_oper_in[24]));

	OBUF QL_INST_F2A_T_22_5 (.IN_OBUF(m0_oper1_rdata_int[23]),.OUT_OBUF(m0_m1_oper_in[23]));

	OBUF QL_INST_F2A_T_22_6 (.IN_OBUF(m0_oper1_rdata_int[22]),.OUT_OBUF(m0_m1_oper_in[22]));

	OBUF QL_INST_F2A_T_22_7 (.IN_OBUF(m0_oper1_rdata_int[21]),.OUT_OBUF(m0_m1_oper_in[21]));

	OBUF QL_INST_F2A_T_22_8 (.IN_OBUF(m0_oper1_rdata_int[20]),.OUT_OBUF(m0_m1_oper_in[20]));

	OBUF QL_INST_F2A_T_22_9 (.IN_OBUF(m0_oper1_rdata_int[19]),.OUT_OBUF(m0_m1_oper_in[19]));

	OBUF QL_INST_F2A_T_22_10 (.IN_OBUF(m0_oper1_rdata_int[18]),.OUT_OBUF(m0_m1_oper_in[18]));

	OBUF QL_INST_F2A_T_22_11 (.IN_OBUF(m0_oper1_rdata_int[17]),.OUT_OBUF(m0_m1_oper_in[17]));

	OBUF QL_INST_F2A_T_22_12 (.IN_OBUF(m0_oper1_rdata_int[16]),.OUT_OBUF(m0_m1_oper_in[16]));

	OBUF QL_INST_F2A_T_22_13 (.IN_OBUF(m0_oper1_rdata_int[15]),.OUT_OBUF(m0_m1_oper_in[15]));

	OBUF QL_INST_F2A_T_22_14 (.IN_OBUF(m0_oper1_rdata_int[14]),.OUT_OBUF(m0_m1_oper_in[14]));

	OBUF QL_INST_F2A_T_22_15 (.IN_OBUF(m0_oper1_rdata_int[13]),.OUT_OBUF(m0_m1_oper_in[13]));

	OBUF QL_INST_F2A_T_22_16 (.IN_OBUF(m0_oper1_rdata_int[12]),.OUT_OBUF(m0_m1_oper_in[12]));

	OBUF QL_INST_F2A_T_22_17 (.IN_OBUF(m0_oper1_rdata_int[11]),.OUT_OBUF(m0_m1_oper_in[11]));

	IBUF QL_INST_A2F_T_22_0 (.IN_IBUF(m0_m1_dataout[4]),.OUT_IBUF(m0_m1_dataout_int[4]));

	IBUF QL_INST_A2F_T_22_1 (.IN_IBUF(m0_m1_dataout[3]),.OUT_IBUF(m0_m1_dataout_int[3]));

	IBUF QL_INST_A2F_T_22_2 (.IN_IBUF(m0_m1_dataout[2]),.OUT_IBUF(m0_m1_dataout_int[2]));

	IBUF QL_INST_A2F_T_22_3 (.IN_IBUF(m0_m1_dataout[1]),.OUT_IBUF(m0_m1_dataout_int[1]));

	IBUF QL_INST_A2F_T_22_4 (.IN_IBUF(m0_m1_dataout[0]),.OUT_IBUF(m0_m1_dataout_int[0]));

	OBUF QL_INST_F2A_T_23_0 (.IN_OBUF(m0_oper1_rdata_int[10]),.OUT_OBUF(m0_m1_oper_in[10]));

	OBUF QL_INST_F2A_T_23_1 (.IN_OBUF(m0_oper1_rdata_int[9]),.OUT_OBUF(m0_m1_oper_in[9]));

	OBUF QL_INST_F2A_T_23_2 (.IN_OBUF(m0_oper1_rdata_int[8]),.OUT_OBUF(m0_m1_oper_in[8]));

	OBUF QL_INST_F2A_T_23_3 (.IN_OBUF(m0_oper1_rdata_int[7]),.OUT_OBUF(m0_m1_oper_in[7]));

	OBUF QL_INST_F2A_T_23_4 (.IN_OBUF(m0_oper1_rdata_int[6]),.OUT_OBUF(m0_m1_oper_in[6]));

	OBUF QL_INST_F2A_T_23_5 (.IN_OBUF(m0_oper1_rdata_int[5]),.OUT_OBUF(m0_m1_oper_in[5]));

	OBUF QL_INST_F2A_T_23_6 (.IN_OBUF(m0_oper1_rdata_int[4]),.OUT_OBUF(m0_m1_oper_in[4]));

	OBUF QL_INST_F2A_T_23_7 (.IN_OBUF(m0_oper1_rdata_int[3]),.OUT_OBUF(m0_m1_oper_in[3]));

	OBUF QL_INST_F2A_T_23_8 (.IN_OBUF(m0_oper1_rdata_int[2]),.OUT_OBUF(m0_m1_oper_in[2]));

	OBUF QL_INST_F2A_T_23_9 (.IN_OBUF(m0_oper1_rdata_int[1]),.OUT_OBUF(m0_m1_oper_in[1]));

	OBUF QL_INST_F2A_T_23_10 (.IN_OBUF(m0_oper1_rdata_int[0]),.OUT_OBUF(m0_m1_oper_in[0]));

	OBUF QL_INST_F2A_T_24_16 (.IN_OBUF(m0_oper1_wdata_dup_0[31]),.OUT_OBUF(m0_oper1_wdata[31]));

	OBUF QL_INST_F2A_T_24_17 (.IN_OBUF(m0_oper1_wdata_dup_0[30]),.OUT_OBUF(m0_oper1_wdata[30]));

	DBUF QL_INST_F2Adef_T_24_0 (.IN_DBUF(GND),.OUT_DBUF(m0_oper1_powerdn));

	OBUF QL_INST_F2A_T_25_0 (.IN_OBUF(m0_oper1_wdata_dup_0[29]),.OUT_OBUF(m0_oper1_wdata[29]));

	OBUF QL_INST_F2A_T_25_1 (.IN_OBUF(m0_oper1_wdata_dup_0[28]),.OUT_OBUF(m0_oper1_wdata[28]));

	OBUF QL_INST_F2A_T_25_2 (.IN_OBUF(m0_oper1_wdata_dup_0[27]),.OUT_OBUF(m0_oper1_wdata[27]));

	OBUF QL_INST_F2A_T_25_3 (.IN_OBUF(m0_oper1_wdata_dup_0[26]),.OUT_OBUF(m0_oper1_wdata[26]));

	OBUF QL_INST_F2A_T_25_4 (.IN_OBUF(m0_oper1_wdata_dup_0[25]),.OUT_OBUF(m0_oper1_wdata[25]));

	OBUF QL_INST_F2A_T_25_5 (.IN_OBUF(m0_oper1_wdata_dup_0[24]),.OUT_OBUF(m0_oper1_wdata[24]));

	OBUF QL_INST_F2A_T_25_6 (.IN_OBUF(m0_oper1_wdata_dup_0[23]),.OUT_OBUF(m0_oper1_wdata[23]));

	OBUF QL_INST_F2A_T_25_7 (.IN_OBUF(m0_oper1_wdata_dup_0[22]),.OUT_OBUF(m0_oper1_wdata[22]));

	OBUF QL_INST_F2A_T_25_8 (.IN_OBUF(m0_oper1_wdata_dup_0[21]),.OUT_OBUF(m0_oper1_wdata[21]));

	OBUF QL_INST_F2A_T_25_9 (.IN_OBUF(m0_oper1_wdata_dup_0[20]),.OUT_OBUF(m0_oper1_wdata[20]));

	OBUF QL_INST_F2A_T_25_10 (.IN_OBUF(m0_oper1_wdata_dup_0[19]),.OUT_OBUF(m0_oper1_wdata[19]));

	OBUF QL_INST_F2A_T_25_11 (.IN_OBUF(m0_oper1_wdata_dup_0[18]),.OUT_OBUF(m0_oper1_wdata[18]));

	IBUF QL_INST_A2F_T_25_1 (.IN_IBUF(m0_oper1_rdata[31]),.OUT_IBUF(m0_oper1_rdata_int[31]));

	IBUF QL_INST_A2F_T_25_2 (.IN_IBUF(m0_oper1_rdata[30]),.OUT_IBUF(m0_oper1_rdata_int[30]));

	IBUF QL_INST_A2F_T_25_3 (.IN_IBUF(m0_oper1_rdata[29]),.OUT_IBUF(m0_oper1_rdata_int[29]));

	IBUF QL_INST_A2F_T_25_4 (.IN_IBUF(m0_oper1_rdata[28]),.OUT_IBUF(m0_oper1_rdata_int[28]));

	IBUF QL_INST_A2F_T_25_5 (.IN_IBUF(m0_oper1_rdata[27]),.OUT_IBUF(m0_oper1_rdata_int[27]));

	OBUF QL_INST_F2A_T_26_0 (.IN_OBUF(m0_oper1_wdata_dup_0[17]),.OUT_OBUF(m0_oper1_wdata[17]));

	OBUF QL_INST_F2A_T_26_1 (.IN_OBUF(m0_oper1_wdata_dup_0[16]),.OUT_OBUF(m0_oper1_wdata[16]));

	OBUF QL_INST_F2A_T_26_2 (.IN_OBUF(m0_oper1_wdata_dup_0[15]),.OUT_OBUF(m0_oper1_wdata[15]));

	OBUF QL_INST_F2A_T_26_3 (.IN_OBUF(m0_oper1_wdata_dup_0[14]),.OUT_OBUF(m0_oper1_wdata[14]));

	OBUF QL_INST_F2A_T_26_4 (.IN_OBUF(m0_oper1_wdata_dup_0[13]),.OUT_OBUF(m0_oper1_wdata[13]));

	OBUF QL_INST_F2A_T_26_5 (.IN_OBUF(m0_oper1_wdata_dup_0[12]),.OUT_OBUF(m0_oper1_wdata[12]));

	OBUF QL_INST_F2A_T_26_6 (.IN_OBUF(m0_oper1_wdata_dup_0[11]),.OUT_OBUF(m0_oper1_wdata[11]));

	OBUF QL_INST_F2A_T_26_7 (.IN_OBUF(m0_oper1_wdata_dup_0[10]),.OUT_OBUF(m0_oper1_wdata[10]));

	OBUF QL_INST_F2A_T_26_8 (.IN_OBUF(m0_oper1_wdata_dup_0[9]),.OUT_OBUF(m0_oper1_wdata[9]));

	OBUF QL_INST_F2A_T_26_9 (.IN_OBUF(m0_oper1_wdata_dup_0[8]),.OUT_OBUF(m0_oper1_wdata[8]));

	OBUF QL_INST_F2A_T_26_10 (.IN_OBUF(m0_oper1_wdata_dup_0[7]),.OUT_OBUF(m0_oper1_wdata[7]));

	OBUF QL_INST_F2A_T_26_11 (.IN_OBUF(m0_oper1_wdata_dup_0[6]),.OUT_OBUF(m0_oper1_wdata[6]));

	OBUF QL_INST_F2A_T_26_12 (.IN_OBUF(m0_oper1_wdata_dup_0[5]),.OUT_OBUF(m0_oper1_wdata[5]));

	OBUF QL_INST_F2A_T_26_13 (.IN_OBUF(m0_oper1_wdata_dup_0[4]),.OUT_OBUF(m0_oper1_wdata[4]));

	OBUF QL_INST_F2A_T_26_14 (.IN_OBUF(m0_oper1_wdata_dup_0[3]),.OUT_OBUF(m0_oper1_wdata[3]));

	OBUF QL_INST_F2A_T_26_15 (.IN_OBUF(m0_oper1_wdata_dup_0[2]),.OUT_OBUF(m0_oper1_wdata[2]));

	OBUF QL_INST_F2A_T_26_16 (.IN_OBUF(m0_oper1_wdata_dup_0[1]),.OUT_OBUF(m0_oper1_wdata[1]));

	OBUF QL_INST_F2A_T_26_17 (.IN_OBUF(m0_oper1_wdata_dup_0[0]),.OUT_OBUF(m0_oper1_wdata[0]));

	IBUF QL_INST_A2F_T_26_0 (.IN_IBUF(m0_oper1_rdata[26]),.OUT_IBUF(m0_oper1_rdata_int[26]));

	IBUF QL_INST_A2F_T_26_1 (.IN_IBUF(m0_oper1_rdata[25]),.OUT_IBUF(m0_oper1_rdata_int[25]));

	IBUF QL_INST_A2F_T_26_2 (.IN_IBUF(m0_oper1_rdata[24]),.OUT_IBUF(m0_oper1_rdata_int[24]));

	IBUF QL_INST_A2F_T_26_3 (.IN_IBUF(m0_oper1_rdata[23]),.OUT_IBUF(m0_oper1_rdata_int[23]));

	IBUF QL_INST_A2F_T_26_4 (.IN_IBUF(m0_oper1_rdata[22]),.OUT_IBUF(m0_oper1_rdata_int[22]));

	IBUF QL_INST_A2F_T_26_5 (.IN_IBUF(m0_oper1_rdata[21]),.OUT_IBUF(m0_oper1_rdata_int[21]));

	IBUF QL_INST_A2F_T_26_6 (.IN_IBUF(m0_oper1_rdata[20]),.OUT_IBUF(m0_oper1_rdata_int[20]));

	IBUF QL_INST_A2F_T_26_7 (.IN_IBUF(m0_oper1_rdata[19]),.OUT_IBUF(m0_oper1_rdata_int[19]));

	OBUF QL_INST_F2A_T_27_0 (.IN_OBUF(m0_oper1_waddr_dup_0[11]),.OUT_OBUF(m0_oper1_waddr[11]));

	OBUF QL_INST_F2A_T_27_1 (.IN_OBUF(m0_oper1_waddr_dup_0[10]),.OUT_OBUF(m0_oper1_waddr[10]));

	OBUF QL_INST_F2A_T_27_2 (.IN_OBUF(m0_oper1_waddr_dup_0[9]),.OUT_OBUF(m0_oper1_waddr[9]));

	OBUF QL_INST_F2A_T_27_3 (.IN_OBUF(m0_oper1_waddr_dup_0[8]),.OUT_OBUF(m0_oper1_waddr[8]));

	OBUF QL_INST_F2A_T_27_4 (.IN_OBUF(m0_oper1_waddr_dup_0[7]),.OUT_OBUF(m0_oper1_waddr[7]));

	OBUF QL_INST_F2A_T_27_5 (.IN_OBUF(m0_oper1_waddr_dup_0[6]),.OUT_OBUF(m0_oper1_waddr[6]));

	OBUF QL_INST_F2A_T_27_6 (.IN_OBUF(m0_oper1_waddr_dup_0[5]),.OUT_OBUF(m0_oper1_waddr[5]));

	OBUF QL_INST_F2A_T_27_7 (.IN_OBUF(m0_oper1_waddr_dup_0[4]),.OUT_OBUF(m0_oper1_waddr[4]));

	OBUF QL_INST_F2A_T_27_8 (.IN_OBUF(m0_oper1_waddr_dup_0[3]),.OUT_OBUF(m0_oper1_waddr[3]));

	OBUF QL_INST_F2A_T_27_9 (.IN_OBUF(m0_oper1_waddr_dup_0[2]),.OUT_OBUF(m0_oper1_waddr[2]));

	OBUF QL_INST_F2A_T_27_10 (.IN_OBUF(m0_oper1_waddr_dup_0[1]),.OUT_OBUF(m0_oper1_waddr[1]));

	OBUF QL_INST_F2A_T_27_11 (.IN_OBUF(m0_oper1_waddr_dup_0[0]),.OUT_OBUF(m0_oper1_waddr[0]));

	IBUF QL_INST_A2F_T_27_0 (.IN_IBUF(m0_oper1_rdata[18]),.OUT_IBUF(m0_oper1_rdata_int[18]));

	IBUF QL_INST_A2F_T_27_1 (.IN_IBUF(m0_oper1_rdata[17]),.OUT_IBUF(m0_oper1_rdata_int[17]));

	IBUF QL_INST_A2F_T_27_2 (.IN_IBUF(m0_oper1_rdata[16]),.OUT_IBUF(m0_oper1_rdata_int[16]));

	IBUF QL_INST_A2F_T_27_3 (.IN_IBUF(m0_oper1_rdata[15]),.OUT_IBUF(m0_oper1_rdata_int[15]));

	IBUF QL_INST_A2F_T_27_4 (.IN_IBUF(m0_oper1_rdata[14]),.OUT_IBUF(m0_oper1_rdata_int[14]));

	IBUF QL_INST_A2F_T_27_5 (.IN_IBUF(m0_oper1_rdata[13]),.OUT_IBUF(m0_oper1_rdata_int[13]));

	OBUF QL_INST_F2A_T_28_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_28_padClk),.OUT_OBUF(m0_oper1_wclk));

	OBUF QL_INST_F2A_T_28_1 (.IN_OBUF(m0_oper1_wmode_dup_0[1]),.OUT_OBUF(m0_oper1_wmode[1]));

	OBUF QL_INST_F2A_T_28_2 (.IN_OBUF(m0_oper1_wmode_dup_0[0]),.OUT_OBUF(m0_oper1_wmode[0]));

	OBUF QL_INST_F2A_T_28_3 (.IN_OBUF(m0_oper1_wdsel_dup_0),.OUT_OBUF(m0_oper1_wdsel));

	OBUF QL_INST_F2A_T_28_4 (.IN_OBUF(m0_oper1_we_dup_0),.OUT_OBUF(m0_oper1_we));

	OBUF QL_INST_F2A_T_28_15 (.IN_OBUF(m0_oper1_rmode_dup_0[1]),.OUT_OBUF(m0_oper1_rmode[1]));

	OBUF QL_INST_F2A_T_28_16 (.IN_OBUF(m0_oper1_rmode_dup_0[0]),.OUT_OBUF(m0_oper1_rmode[0]));

	OBUF QL_INST_F2A_T_28_17 (.IN_OBUF(m0_oper1_raddr_dup_0[11]),.OUT_OBUF(m0_oper1_raddr[11]));

	IBUF QL_INST_A2F_T_28_1 (.IN_IBUF(m0_oper1_rdata[12]),.OUT_IBUF(m0_oper1_rdata_int[12]));

	IBUF QL_INST_A2F_T_28_2 (.IN_IBUF(m0_oper1_rdata[11]),.OUT_IBUF(m0_oper1_rdata_int[11]));

	IBUF QL_INST_A2F_T_28_3 (.IN_IBUF(m0_oper1_rdata[10]),.OUT_IBUF(m0_oper1_rdata_int[10]));

	IBUF QL_INST_A2F_T_28_4 (.IN_IBUF(m0_oper1_rdata[9]),.OUT_IBUF(m0_oper1_rdata_int[9]));

	IBUF QL_INST_A2F_T_28_5 (.IN_IBUF(m0_oper1_rdata[8]),.OUT_IBUF(m0_oper1_rdata_int[8]));

	IBUF QL_INST_A2F_T_28_6 (.IN_IBUF(m0_oper1_rdata[7]),.OUT_IBUF(m0_oper1_rdata_int[7]));

	IBUF QL_INST_A2F_T_28_7 (.IN_IBUF(m0_oper1_rdata[6]),.OUT_IBUF(m0_oper1_rdata_int[6]));

	OBUF QL_INST_F2A_T_29_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_29_padClk),.OUT_OBUF(m0_oper1_rclk));

	OBUF QL_INST_F2A_T_29_1 (.IN_OBUF(m0_oper1_raddr_dup_0[10]),.OUT_OBUF(m0_oper1_raddr[10]));

	OBUF QL_INST_F2A_T_29_2 (.IN_OBUF(m0_oper1_raddr_dup_0[9]),.OUT_OBUF(m0_oper1_raddr[9]));

	OBUF QL_INST_F2A_T_29_3 (.IN_OBUF(m0_oper1_raddr_dup_0[8]),.OUT_OBUF(m0_oper1_raddr[8]));

	OBUF QL_INST_F2A_T_29_4 (.IN_OBUF(m0_oper1_raddr_dup_0[7]),.OUT_OBUF(m0_oper1_raddr[7]));

	OBUF QL_INST_F2A_T_29_5 (.IN_OBUF(m0_oper1_raddr_dup_0[6]),.OUT_OBUF(m0_oper1_raddr[6]));

	OBUF QL_INST_F2A_T_29_6 (.IN_OBUF(m0_oper1_raddr_dup_0[5]),.OUT_OBUF(m0_oper1_raddr[5]));

	OBUF QL_INST_F2A_T_29_7 (.IN_OBUF(m0_oper1_raddr_dup_0[4]),.OUT_OBUF(m0_oper1_raddr[4]));

	OBUF QL_INST_F2A_T_29_8 (.IN_OBUF(m0_oper1_raddr_dup_0[3]),.OUT_OBUF(m0_oper1_raddr[3]));

	OBUF QL_INST_F2A_T_29_9 (.IN_OBUF(m0_oper1_raddr_dup_0[2]),.OUT_OBUF(m0_oper1_raddr[2]));

	OBUF QL_INST_F2A_T_29_10 (.IN_OBUF(m0_oper1_raddr_dup_0[1]),.OUT_OBUF(m0_oper1_raddr[1]));

	OBUF QL_INST_F2A_T_29_11 (.IN_OBUF(m0_oper1_raddr_dup_0[0]),.OUT_OBUF(m0_oper1_raddr[0]));

	IBUF QL_INST_A2F_T_29_0 (.IN_IBUF(m0_oper1_rdata[5]),.OUT_IBUF(m0_oper1_rdata_int[5]));

	IBUF QL_INST_A2F_T_29_1 (.IN_IBUF(m0_oper1_rdata[4]),.OUT_IBUF(m0_oper1_rdata_int[4]));

	IBUF QL_INST_A2F_T_29_2 (.IN_IBUF(m0_oper1_rdata[3]),.OUT_IBUF(m0_oper1_rdata_int[3]));

	IBUF QL_INST_A2F_T_29_3 (.IN_IBUF(m0_oper1_rdata[2]),.OUT_IBUF(m0_oper1_rdata_int[2]));

	IBUF QL_INST_A2F_T_29_4 (.IN_IBUF(m0_oper1_rdata[1]),.OUT_IBUF(m0_oper1_rdata_int[1]));

	IBUF QL_INST_A2F_T_29_5 (.IN_IBUF(m0_oper1_rdata[0]),.OUT_IBUF(m0_oper1_rdata_int[0]));

	OBUF QL_INST_F2A_R_3_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_33_padClk),.OUT_OBUF(tcdm_clk_p0));

	OBUF QL_INST_F2A_R_3_1 (.IN_OBUF(tcdm_req_p0_dup_0),.OUT_OBUF(tcdm_req_p0));

	OBUF QL_INST_F2A_R_3_2 (.IN_OBUF(tcdm_wen_p0_dup_0),.OUT_OBUF(tcdm_wen_p0));

	OBUF QL_INST_F2A_R_3_3 (.IN_OBUF(tcdm_be_p0_dup_0[0]),.OUT_OBUF(tcdm_be_p0[0]));

	OBUF QL_INST_F2A_R_3_4 (.IN_OBUF(tcdm_be_p0_dup_0[1]),.OUT_OBUF(tcdm_be_p0[1]));

	OBUF QL_INST_F2A_R_3_5 (.IN_OBUF(tcdm_be_p0_dup_0[2]),.OUT_OBUF(tcdm_be_p0[2]));

	OBUF QL_INST_F2A_R_3_6 (.IN_OBUF(tcdm_be_p0_dup_0[3]),.OUT_OBUF(tcdm_be_p0[3]));

	OBUF QL_INST_F2A_R_3_8 (.IN_OBUF(tcdm_addr_p0_dup_0[0]),.OUT_OBUF(tcdm_addr_p0[0]));

	OBUF QL_INST_F2A_R_3_9 (.IN_OBUF(tcdm_addr_p0_dup_0[1]),.OUT_OBUF(tcdm_addr_p0[1]));

	OBUF QL_INST_F2A_R_3_10 (.IN_OBUF(tcdm_addr_p0_dup_0[2]),.OUT_OBUF(tcdm_addr_p0[2]));

	OBUF QL_INST_F2A_R_3_11 (.IN_OBUF(tcdm_addr_p0_dup_0[3]),.OUT_OBUF(tcdm_addr_p0[3]));

	IBUF QL_INST_A2F_R_3_0 (.IN_IBUF(tcdm_rdata_p0[0]),.OUT_IBUF(tcdm_rdata_p0_int[0]));

	IBUF QL_INST_A2F_R_3_1 (.IN_IBUF(tcdm_rdata_p0[1]),.OUT_IBUF(tcdm_rdata_p0_int[1]));

	IBUF QL_INST_A2F_R_3_2 (.IN_IBUF(tcdm_rdata_p0[2]),.OUT_IBUF(tcdm_rdata_p0_int[2]));

	IBUF QL_INST_A2F_R_3_3 (.IN_IBUF(tcdm_rdata_p0[3]),.OUT_IBUF(tcdm_rdata_p0_int[3]));

	IBUF QL_INST_A2F_R_3_4 (.IN_IBUF(tcdm_valid_p0),.OUT_IBUF(tcdm_valid_p0_int));

	IBUF QL_INST_A2F_R_3_5 (.IN_IBUF(tcdm_gnt_p0),.OUT_IBUF(tcdm_gnt_p0_int));

	OBUF QL_INST_F2A_R_4_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[0]),.OUT_OBUF(tcdm_wdata_p0[0]));

	OBUF QL_INST_F2A_R_4_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[1]),.OUT_OBUF(tcdm_wdata_p0[1]));

	OBUF QL_INST_F2A_R_4_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[2]),.OUT_OBUF(tcdm_wdata_p0[2]));

	OBUF QL_INST_F2A_R_4_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[3]),.OUT_OBUF(tcdm_wdata_p0[3]));

	OBUF QL_INST_F2A_R_4_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[4]),.OUT_OBUF(tcdm_wdata_p0[4]));

	OBUF QL_INST_F2A_R_4_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[5]),.OUT_OBUF(tcdm_wdata_p0[5]));

	OBUF QL_INST_F2A_R_4_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[6]),.OUT_OBUF(tcdm_wdata_p0[6]));

	OBUF QL_INST_F2A_R_4_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[7]),.OUT_OBUF(tcdm_wdata_p0[7]));

	OBUF QL_INST_F2A_R_4_9 (.IN_OBUF(tcdm_addr_p0_dup_0[4]),.OUT_OBUF(tcdm_addr_p0[4]));

	OBUF QL_INST_F2A_R_4_10 (.IN_OBUF(tcdm_addr_p0_dup_0[5]),.OUT_OBUF(tcdm_addr_p0[5]));

	OBUF QL_INST_F2A_R_4_11 (.IN_OBUF(tcdm_addr_p0_dup_0[6]),.OUT_OBUF(tcdm_addr_p0[6]));

	OBUF QL_INST_F2A_R_4_12 (.IN_OBUF(tcdm_addr_p0_dup_0[7]),.OUT_OBUF(tcdm_addr_p0[7]));

	OBUF QL_INST_F2A_R_4_13 (.IN_OBUF(tcdm_addr_p0_dup_0[8]),.OUT_OBUF(tcdm_addr_p0[8]));

	OBUF QL_INST_F2A_R_4_14 (.IN_OBUF(tcdm_addr_p0_dup_0[9]),.OUT_OBUF(tcdm_addr_p0[9]));

	IBUF QL_INST_A2F_R_4_0 (.IN_IBUF(tcdm_rdata_p0[4]),.OUT_IBUF(tcdm_rdata_p0_int[4]));

	IBUF QL_INST_A2F_R_4_1 (.IN_IBUF(tcdm_rdata_p0[5]),.OUT_IBUF(tcdm_rdata_p0_int[5]));

	IBUF QL_INST_A2F_R_4_2 (.IN_IBUF(tcdm_rdata_p0[6]),.OUT_IBUF(tcdm_rdata_p0_int[6]));

	IBUF QL_INST_A2F_R_4_3 (.IN_IBUF(tcdm_rdata_p0[7]),.OUT_IBUF(tcdm_rdata_p0_int[7]));

	IBUF QL_INST_A2F_R_4_4 (.IN_IBUF(tcdm_rdata_p0[8]),.OUT_IBUF(tcdm_rdata_p0_int[8]));

	IBUF QL_INST_A2F_R_4_5 (.IN_IBUF(tcdm_rdata_p0[9]),.OUT_IBUF(tcdm_rdata_p0_int[9]));

	IBUF QL_INST_A2F_R_4_6 (.IN_IBUF(tcdm_rdata_p0[10]),.OUT_IBUF(tcdm_rdata_p0_int[10]));

	IBUF QL_INST_A2F_R_4_7 (.IN_IBUF(tcdm_rdata_p0[11]),.OUT_IBUF(tcdm_rdata_p0_int[11]));

	OBUF QL_INST_F2A_R_5_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[8]),.OUT_OBUF(tcdm_wdata_p0[8]));

	OBUF QL_INST_F2A_R_5_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[9]),.OUT_OBUF(tcdm_wdata_p0[9]));

	OBUF QL_INST_F2A_R_5_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[10]),.OUT_OBUF(tcdm_wdata_p0[10]));

	OBUF QL_INST_F2A_R_5_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[11]),.OUT_OBUF(tcdm_wdata_p0[11]));

	OBUF QL_INST_F2A_R_5_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[12]),.OUT_OBUF(tcdm_wdata_p0[12]));

	OBUF QL_INST_F2A_R_5_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[13]),.OUT_OBUF(tcdm_wdata_p0[13]));

	OBUF QL_INST_F2A_R_5_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[14]),.OUT_OBUF(tcdm_wdata_p0[14]));

	OBUF QL_INST_F2A_R_5_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[15]),.OUT_OBUF(tcdm_wdata_p0[15]));

	OBUF QL_INST_F2A_R_5_8 (.IN_OBUF(tcdm_addr_p0_dup_0[10]),.OUT_OBUF(tcdm_addr_p0[10]));

	OBUF QL_INST_F2A_R_5_9 (.IN_OBUF(tcdm_addr_p0_dup_0[11]),.OUT_OBUF(tcdm_addr_p0[11]));

	OBUF QL_INST_F2A_R_5_10 (.IN_OBUF(tcdm_addr_p0_dup_0[12]),.OUT_OBUF(tcdm_addr_p0[12]));

	OBUF QL_INST_F2A_R_5_11 (.IN_OBUF(tcdm_addr_p0_dup_0[13]),.OUT_OBUF(tcdm_addr_p0[13]));

	IBUF QL_INST_A2F_R_5_0 (.IN_IBUF(tcdm_rdata_p0[12]),.OUT_IBUF(tcdm_rdata_p0_int[12]));

	IBUF QL_INST_A2F_R_5_1 (.IN_IBUF(tcdm_rdata_p0[13]),.OUT_IBUF(tcdm_rdata_p0_int[13]));

	IBUF QL_INST_A2F_R_5_2 (.IN_IBUF(tcdm_rdata_p0[14]),.OUT_IBUF(tcdm_rdata_p0_int[14]));

	IBUF QL_INST_A2F_R_5_3 (.IN_IBUF(tcdm_rdata_p0[15]),.OUT_IBUF(tcdm_rdata_p0_int[15]));

	OBUF QL_INST_F2A_R_6_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[16]),.OUT_OBUF(tcdm_wdata_p0[16]));

	OBUF QL_INST_F2A_R_6_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[17]),.OUT_OBUF(tcdm_wdata_p0[17]));

	OBUF QL_INST_F2A_R_6_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[18]),.OUT_OBUF(tcdm_wdata_p0[18]));

	OBUF QL_INST_F2A_R_6_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[19]),.OUT_OBUF(tcdm_wdata_p0[19]));

	OBUF QL_INST_F2A_R_6_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[20]),.OUT_OBUF(tcdm_wdata_p0[20]));

	OBUF QL_INST_F2A_R_6_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[21]),.OUT_OBUF(tcdm_wdata_p0[21]));

	OBUF QL_INST_F2A_R_6_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[22]),.OUT_OBUF(tcdm_wdata_p0[22]));

	OBUF QL_INST_F2A_R_6_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[23]),.OUT_OBUF(tcdm_wdata_p0[23]));

	OBUF QL_INST_F2A_R_6_12 (.IN_OBUF(tcdm_addr_p0_dup_0[14]),.OUT_OBUF(tcdm_addr_p0[14]));

	OBUF QL_INST_F2A_R_6_13 (.IN_OBUF(tcdm_addr_p0_dup_0[15]),.OUT_OBUF(tcdm_addr_p0[15]));

	OBUF QL_INST_F2A_R_6_14 (.IN_OBUF(tcdm_addr_p0_dup_0[16]),.OUT_OBUF(tcdm_addr_p0[16]));

	OBUF QL_INST_F2A_R_6_15 (.IN_OBUF(tcdm_addr_p0_dup_0[17]),.OUT_OBUF(tcdm_addr_p0[17]));

	OBUF QL_INST_F2A_R_6_16 (.IN_OBUF(tcdm_addr_p0_dup_0[18]),.OUT_OBUF(tcdm_addr_p0[18]));

	OBUF QL_INST_F2A_R_6_17 (.IN_OBUF(tcdm_addr_p0_dup_0[19]),.OUT_OBUF(tcdm_addr_p0[19]));

	IBUF QL_INST_A2F_R_6_0 (.IN_IBUF(RESET[0]),.OUT_IBUF(RESET_int[0]));

	IBUF QL_INST_A2F_R_6_1 (.IN_IBUF(tcdm_rdata_p0[16]),.OUT_IBUF(tcdm_rdata_p0_int[16]));

	IBUF QL_INST_A2F_R_6_2 (.IN_IBUF(tcdm_rdata_p0[17]),.OUT_IBUF(tcdm_rdata_p0_int[17]));

	IBUF QL_INST_A2F_R_6_3 (.IN_IBUF(tcdm_rdata_p0[18]),.OUT_IBUF(tcdm_rdata_p0_int[18]));

	IBUF QL_INST_A2F_R_6_4 (.IN_IBUF(tcdm_rdata_p0[19]),.OUT_IBUF(tcdm_rdata_p0_int[19]));

	IBUF QL_INST_A2F_R_6_5 (.IN_IBUF(tcdm_rdata_p0[20]),.OUT_IBUF(tcdm_rdata_p0_int[20]));

	IBUF QL_INST_A2F_R_6_6 (.IN_IBUF(tcdm_rdata_p0[21]),.OUT_IBUF(tcdm_rdata_p0_int[21]));

	OBUF QL_INST_F2A_R_7_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[24]),.OUT_OBUF(tcdm_wdata_p0[24]));

	OBUF QL_INST_F2A_R_7_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[25]),.OUT_OBUF(tcdm_wdata_p0[25]));

	OBUF QL_INST_F2A_R_7_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[26]),.OUT_OBUF(tcdm_wdata_p0[26]));

	OBUF QL_INST_F2A_R_7_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[27]),.OUT_OBUF(tcdm_wdata_p0[27]));

	OBUF QL_INST_F2A_R_7_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[28]),.OUT_OBUF(tcdm_wdata_p0[28]));

	OBUF QL_INST_F2A_R_7_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[29]),.OUT_OBUF(tcdm_wdata_p0[29]));

	OBUF QL_INST_F2A_R_7_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[30]),.OUT_OBUF(tcdm_wdata_p0[30]));

	OBUF QL_INST_F2A_R_7_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[31]),.OUT_OBUF(tcdm_wdata_p0[31]));

	IBUF QL_INST_A2F_R_7_0 (.IN_IBUF(tcdm_rdata_p0[22]),.OUT_IBUF(tcdm_rdata_p0_int[22]));

	IBUF QL_INST_A2F_R_7_1 (.IN_IBUF(tcdm_rdata_p0[23]),.OUT_IBUF(tcdm_rdata_p0_int[23]));

	IBUF QL_INST_A2F_R_7_2 (.IN_IBUF(tcdm_rdata_p0[24]),.OUT_IBUF(tcdm_rdata_p0_int[24]));

	IBUF QL_INST_A2F_R_7_3 (.IN_IBUF(tcdm_rdata_p0[25]),.OUT_IBUF(tcdm_rdata_p0_int[25]));

	IBUF QL_INST_A2F_R_7_4 (.IN_IBUF(tcdm_rdata_p0[26]),.OUT_IBUF(tcdm_rdata_p0_int[26]));

	IBUF QL_INST_A2F_R_7_5 (.IN_IBUF(tcdm_rdata_p0[27]),.OUT_IBUF(tcdm_rdata_p0_int[27]));

	IBUF QL_INST_A2F_R_8_0 (.IN_IBUF(tcdm_rdata_p0[28]),.OUT_IBUF(tcdm_rdata_p0_int[28]));

	IBUF QL_INST_A2F_R_8_1 (.IN_IBUF(tcdm_rdata_p0[29]),.OUT_IBUF(tcdm_rdata_p0_int[29]));

	IBUF QL_INST_A2F_R_8_2 (.IN_IBUF(tcdm_rdata_p0[30]),.OUT_IBUF(tcdm_rdata_p0_int[30]));

	IBUF QL_INST_A2F_R_8_3 (.IN_IBUF(tcdm_rdata_p0[31]),.OUT_IBUF(tcdm_rdata_p0_int[31]));

	OBUF QL_INST_F2A_R_9_0 (.IN_OBUF(CLK_int_0__CAND0_TRSBR_33_padClk),.OUT_OBUF(tcdm_clk_p1));

	OBUF QL_INST_F2A_R_9_1 (.IN_OBUF(tcdm_req_p1_dup_0),.OUT_OBUF(tcdm_req_p1));

	OBUF QL_INST_F2A_R_9_2 (.IN_OBUF(tcdm_wen_p1_dup_0),.OUT_OBUF(tcdm_wen_p1));

	OBUF QL_INST_F2A_R_9_3 (.IN_OBUF(tcdm_be_p1_dup_0[0]),.OUT_OBUF(tcdm_be_p1[0]));

	OBUF QL_INST_F2A_R_9_4 (.IN_OBUF(tcdm_be_p1_dup_0[1]),.OUT_OBUF(tcdm_be_p1[1]));

	OBUF QL_INST_F2A_R_9_5 (.IN_OBUF(tcdm_be_p1_dup_0[2]),.OUT_OBUF(tcdm_be_p1[2]));

	OBUF QL_INST_F2A_R_9_6 (.IN_OBUF(tcdm_be_p1_dup_0[3]),.OUT_OBUF(tcdm_be_p1[3]));

	OBUF QL_INST_F2A_R_9_8 (.IN_OBUF(tcdm_addr_p1_dup_0[0]),.OUT_OBUF(tcdm_addr_p1[0]));

	OBUF QL_INST_F2A_R_9_9 (.IN_OBUF(tcdm_addr_p1_dup_0[1]),.OUT_OBUF(tcdm_addr_p1[1]));

	OBUF QL_INST_F2A_R_9_10 (.IN_OBUF(tcdm_addr_p1_dup_0[2]),.OUT_OBUF(tcdm_addr_p1[2]));

	OBUF QL_INST_F2A_R_9_11 (.IN_OBUF(tcdm_addr_p1_dup_0[3]),.OUT_OBUF(tcdm_addr_p1[3]));

	IBUF QL_INST_A2F_R_9_0 (.IN_IBUF(tcdm_rdata_p1[0]),.OUT_IBUF(tcdm_rdata_p1_int[0]));

	IBUF QL_INST_A2F_R_9_1 (.IN_IBUF(tcdm_rdata_p1[1]),.OUT_IBUF(tcdm_rdata_p1_int[1]));

	IBUF QL_INST_A2F_R_9_2 (.IN_IBUF(tcdm_rdata_p1[2]),.OUT_IBUF(tcdm_rdata_p1_int[2]));

	IBUF QL_INST_A2F_R_9_3 (.IN_IBUF(tcdm_rdata_p1[3]),.OUT_IBUF(tcdm_rdata_p1_int[3]));

	IBUF QL_INST_A2F_R_9_4 (.IN_IBUF(tcdm_valid_p1),.OUT_IBUF(tcdm_valid_p1_int));

	IBUF QL_INST_A2F_R_9_5 (.IN_IBUF(tcdm_gnt_p1),.OUT_IBUF(tcdm_gnt_p1_int));

	OBUF QL_INST_F2A_R_10_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[0]),.OUT_OBUF(tcdm_wdata_p1[0]));

	OBUF QL_INST_F2A_R_10_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[1]),.OUT_OBUF(tcdm_wdata_p1[1]));

	OBUF QL_INST_F2A_R_10_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[2]),.OUT_OBUF(tcdm_wdata_p1[2]));

	OBUF QL_INST_F2A_R_10_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[3]),.OUT_OBUF(tcdm_wdata_p1[3]));

	OBUF QL_INST_F2A_R_10_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[4]),.OUT_OBUF(tcdm_wdata_p1[4]));

	OBUF QL_INST_F2A_R_10_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[5]),.OUT_OBUF(tcdm_wdata_p1[5]));

	OBUF QL_INST_F2A_R_10_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[6]),.OUT_OBUF(tcdm_wdata_p1[6]));

	OBUF QL_INST_F2A_R_10_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[7]),.OUT_OBUF(tcdm_wdata_p1[7]));

	OBUF QL_INST_F2A_R_10_9 (.IN_OBUF(tcdm_addr_p1_dup_0[4]),.OUT_OBUF(tcdm_addr_p1[4]));

	OBUF QL_INST_F2A_R_10_10 (.IN_OBUF(tcdm_addr_p1_dup_0[5]),.OUT_OBUF(tcdm_addr_p1[5]));

	OBUF QL_INST_F2A_R_10_11 (.IN_OBUF(tcdm_addr_p1_dup_0[6]),.OUT_OBUF(tcdm_addr_p1[6]));

	OBUF QL_INST_F2A_R_10_12 (.IN_OBUF(tcdm_addr_p1_dup_0[7]),.OUT_OBUF(tcdm_addr_p1[7]));

	OBUF QL_INST_F2A_R_10_13 (.IN_OBUF(tcdm_addr_p1_dup_0[8]),.OUT_OBUF(tcdm_addr_p1[8]));

	OBUF QL_INST_F2A_R_10_14 (.IN_OBUF(tcdm_addr_p1_dup_0[9]),.OUT_OBUF(tcdm_addr_p1[9]));

	IBUF QL_INST_A2F_R_10_0 (.IN_IBUF(tcdm_rdata_p1[4]),.OUT_IBUF(tcdm_rdata_p1_int[4]));

	IBUF QL_INST_A2F_R_10_1 (.IN_IBUF(tcdm_rdata_p1[5]),.OUT_IBUF(tcdm_rdata_p1_int[5]));

	IBUF QL_INST_A2F_R_10_2 (.IN_IBUF(tcdm_rdata_p1[6]),.OUT_IBUF(tcdm_rdata_p1_int[6]));

	IBUF QL_INST_A2F_R_10_3 (.IN_IBUF(tcdm_rdata_p1[7]),.OUT_IBUF(tcdm_rdata_p1_int[7]));

	IBUF QL_INST_A2F_R_10_4 (.IN_IBUF(tcdm_rdata_p1[8]),.OUT_IBUF(tcdm_rdata_p1_int[8]));

	IBUF QL_INST_A2F_R_10_5 (.IN_IBUF(tcdm_rdata_p1[9]),.OUT_IBUF(tcdm_rdata_p1_int[9]));

	IBUF QL_INST_A2F_R_10_6 (.IN_IBUF(tcdm_rdata_p1[10]),.OUT_IBUF(tcdm_rdata_p1_int[10]));

	IBUF QL_INST_A2F_R_10_7 (.IN_IBUF(tcdm_rdata_p1[11]),.OUT_IBUF(tcdm_rdata_p1_int[11]));

	OBUF QL_INST_F2A_R_11_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[8]),.OUT_OBUF(tcdm_wdata_p1[8]));

	OBUF QL_INST_F2A_R_11_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[9]),.OUT_OBUF(tcdm_wdata_p1[9]));

	OBUF QL_INST_F2A_R_11_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[10]),.OUT_OBUF(tcdm_wdata_p1[10]));

	OBUF QL_INST_F2A_R_11_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[11]),.OUT_OBUF(tcdm_wdata_p1[11]));

	OBUF QL_INST_F2A_R_11_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[12]),.OUT_OBUF(tcdm_wdata_p1[12]));

	OBUF QL_INST_F2A_R_11_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[13]),.OUT_OBUF(tcdm_wdata_p1[13]));

	OBUF QL_INST_F2A_R_11_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[14]),.OUT_OBUF(tcdm_wdata_p1[14]));

	OBUF QL_INST_F2A_R_11_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[15]),.OUT_OBUF(tcdm_wdata_p1[15]));

	OBUF QL_INST_F2A_R_11_8 (.IN_OBUF(tcdm_addr_p1_dup_0[10]),.OUT_OBUF(tcdm_addr_p1[10]));

	OBUF QL_INST_F2A_R_11_9 (.IN_OBUF(tcdm_addr_p1_dup_0[11]),.OUT_OBUF(tcdm_addr_p1[11]));

	OBUF QL_INST_F2A_R_11_10 (.IN_OBUF(tcdm_addr_p1_dup_0[12]),.OUT_OBUF(tcdm_addr_p1[12]));

	OBUF QL_INST_F2A_R_11_11 (.IN_OBUF(tcdm_addr_p1_dup_0[13]),.OUT_OBUF(tcdm_addr_p1[13]));

	IBUF QL_INST_A2F_R_11_0 (.IN_IBUF(tcdm_rdata_p1[12]),.OUT_IBUF(tcdm_rdata_p1_int[12]));

	IBUF QL_INST_A2F_R_11_1 (.IN_IBUF(tcdm_rdata_p1[13]),.OUT_IBUF(tcdm_rdata_p1_int[13]));

	IBUF QL_INST_A2F_R_11_2 (.IN_IBUF(tcdm_rdata_p1[14]),.OUT_IBUF(tcdm_rdata_p1_int[14]));

	IBUF QL_INST_A2F_R_11_3 (.IN_IBUF(tcdm_rdata_p1[15]),.OUT_IBUF(tcdm_rdata_p1_int[15]));

	OBUF QL_INST_F2A_R_12_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[16]),.OUT_OBUF(tcdm_wdata_p1[16]));

	OBUF QL_INST_F2A_R_12_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[17]),.OUT_OBUF(tcdm_wdata_p1[17]));

	OBUF QL_INST_F2A_R_12_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[18]),.OUT_OBUF(tcdm_wdata_p1[18]));

	OBUF QL_INST_F2A_R_12_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[19]),.OUT_OBUF(tcdm_wdata_p1[19]));

	OBUF QL_INST_F2A_R_12_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[20]),.OUT_OBUF(tcdm_wdata_p1[20]));

	OBUF QL_INST_F2A_R_12_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[21]),.OUT_OBUF(tcdm_wdata_p1[21]));

	OBUF QL_INST_F2A_R_12_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[22]),.OUT_OBUF(tcdm_wdata_p1[22]));

	OBUF QL_INST_F2A_R_12_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[23]),.OUT_OBUF(tcdm_wdata_p1[23]));

	OBUF QL_INST_F2A_R_12_12 (.IN_OBUF(tcdm_addr_p1_dup_0[14]),.OUT_OBUF(tcdm_addr_p1[14]));

	OBUF QL_INST_F2A_R_12_13 (.IN_OBUF(tcdm_addr_p1_dup_0[15]),.OUT_OBUF(tcdm_addr_p1[15]));

	OBUF QL_INST_F2A_R_12_14 (.IN_OBUF(tcdm_addr_p1_dup_0[16]),.OUT_OBUF(tcdm_addr_p1[16]));

	OBUF QL_INST_F2A_R_12_15 (.IN_OBUF(tcdm_addr_p1_dup_0[17]),.OUT_OBUF(tcdm_addr_p1[17]));

	OBUF QL_INST_F2A_R_12_16 (.IN_OBUF(tcdm_addr_p1_dup_0[18]),.OUT_OBUF(tcdm_addr_p1[18]));

	OBUF QL_INST_F2A_R_12_17 (.IN_OBUF(tcdm_addr_p1_dup_0[19]),.OUT_OBUF(tcdm_addr_p1[19]));

	IBUF QL_INST_A2F_R_12_1 (.IN_IBUF(tcdm_rdata_p1[16]),.OUT_IBUF(tcdm_rdata_p1_int[16]));

	IBUF QL_INST_A2F_R_12_2 (.IN_IBUF(tcdm_rdata_p1[17]),.OUT_IBUF(tcdm_rdata_p1_int[17]));

	IBUF QL_INST_A2F_R_12_3 (.IN_IBUF(tcdm_rdata_p1[18]),.OUT_IBUF(tcdm_rdata_p1_int[18]));

	IBUF QL_INST_A2F_R_12_4 (.IN_IBUF(tcdm_rdata_p1[19]),.OUT_IBUF(tcdm_rdata_p1_int[19]));

	IBUF QL_INST_A2F_R_12_5 (.IN_IBUF(tcdm_rdata_p1[20]),.OUT_IBUF(tcdm_rdata_p1_int[20]));

	IBUF QL_INST_A2F_R_12_6 (.IN_IBUF(tcdm_rdata_p1[21]),.OUT_IBUF(tcdm_rdata_p1_int[21]));

	OBUF QL_INST_F2A_R_13_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[24]),.OUT_OBUF(tcdm_wdata_p1[24]));

	OBUF QL_INST_F2A_R_13_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[25]),.OUT_OBUF(tcdm_wdata_p1[25]));

	OBUF QL_INST_F2A_R_13_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[26]),.OUT_OBUF(tcdm_wdata_p1[26]));

	OBUF QL_INST_F2A_R_13_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[27]),.OUT_OBUF(tcdm_wdata_p1[27]));

	OBUF QL_INST_F2A_R_13_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[28]),.OUT_OBUF(tcdm_wdata_p1[28]));

	OBUF QL_INST_F2A_R_13_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[29]),.OUT_OBUF(tcdm_wdata_p1[29]));

	OBUF QL_INST_F2A_R_13_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[30]),.OUT_OBUF(tcdm_wdata_p1[30]));

	OBUF QL_INST_F2A_R_13_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[31]),.OUT_OBUF(tcdm_wdata_p1[31]));

	IBUF QL_INST_A2F_R_13_0 (.IN_IBUF(tcdm_rdata_p1[22]),.OUT_IBUF(tcdm_rdata_p1_int[22]));

	IBUF QL_INST_A2F_R_13_1 (.IN_IBUF(tcdm_rdata_p1[23]),.OUT_IBUF(tcdm_rdata_p1_int[23]));

	IBUF QL_INST_A2F_R_13_2 (.IN_IBUF(tcdm_rdata_p1[24]),.OUT_IBUF(tcdm_rdata_p1_int[24]));

	IBUF QL_INST_A2F_R_13_3 (.IN_IBUF(tcdm_rdata_p1[25]),.OUT_IBUF(tcdm_rdata_p1_int[25]));

	IBUF QL_INST_A2F_R_13_4 (.IN_IBUF(tcdm_rdata_p1[26]),.OUT_IBUF(tcdm_rdata_p1_int[26]));

	IBUF QL_INST_A2F_R_13_5 (.IN_IBUF(tcdm_rdata_p1[27]),.OUT_IBUF(tcdm_rdata_p1_int[27]));

	IBUF QL_INST_A2F_R_14_0 (.IN_IBUF(tcdm_rdata_p1[28]),.OUT_IBUF(tcdm_rdata_p1_int[28]));

	IBUF QL_INST_A2F_R_14_1 (.IN_IBUF(tcdm_rdata_p1[29]),.OUT_IBUF(tcdm_rdata_p1_int[29]));

	IBUF QL_INST_A2F_R_14_2 (.IN_IBUF(tcdm_rdata_p1[30]),.OUT_IBUF(tcdm_rdata_p1_int[30]));

	IBUF QL_INST_A2F_R_14_3 (.IN_IBUF(tcdm_rdata_p1[31]),.OUT_IBUF(tcdm_rdata_p1_int[31]));

	OBUF QL_INST_F2A_R_17_0 (.IN_OBUF(CLK_int_0__CAND0_BRSTR_33_padClk),.OUT_OBUF(tcdm_clk_p2));

	OBUF QL_INST_F2A_R_17_1 (.IN_OBUF(tcdm_req_p2_dup_0),.OUT_OBUF(tcdm_req_p2));

	OBUF QL_INST_F2A_R_17_2 (.IN_OBUF(tcdm_wen_p2_dup_0),.OUT_OBUF(tcdm_wen_p2));

	OBUF QL_INST_F2A_R_17_3 (.IN_OBUF(tcdm_be_p2_dup_0[0]),.OUT_OBUF(tcdm_be_p2[0]));

	OBUF QL_INST_F2A_R_17_4 (.IN_OBUF(tcdm_be_p2_dup_0[1]),.OUT_OBUF(tcdm_be_p2[1]));

	OBUF QL_INST_F2A_R_17_5 (.IN_OBUF(tcdm_be_p2_dup_0[2]),.OUT_OBUF(tcdm_be_p2[2]));

	OBUF QL_INST_F2A_R_17_6 (.IN_OBUF(tcdm_be_p2_dup_0[3]),.OUT_OBUF(tcdm_be_p2[3]));

	OBUF QL_INST_F2A_R_17_8 (.IN_OBUF(tcdm_addr_p2_dup_0[0]),.OUT_OBUF(tcdm_addr_p2[0]));

	OBUF QL_INST_F2A_R_17_9 (.IN_OBUF(tcdm_addr_p2_dup_0[1]),.OUT_OBUF(tcdm_addr_p2[1]));

	OBUF QL_INST_F2A_R_17_10 (.IN_OBUF(tcdm_addr_p2_dup_0[2]),.OUT_OBUF(tcdm_addr_p2[2]));

	OBUF QL_INST_F2A_R_17_11 (.IN_OBUF(tcdm_addr_p2_dup_0[3]),.OUT_OBUF(tcdm_addr_p2[3]));

	IBUF QL_INST_A2F_R_17_0 (.IN_IBUF(tcdm_rdata_p2[0]),.OUT_IBUF(tcdm_rdata_p2_int[0]));

	IBUF QL_INST_A2F_R_17_1 (.IN_IBUF(tcdm_rdata_p2[1]),.OUT_IBUF(tcdm_rdata_p2_int[1]));

	IBUF QL_INST_A2F_R_17_2 (.IN_IBUF(tcdm_rdata_p2[2]),.OUT_IBUF(tcdm_rdata_p2_int[2]));

	IBUF QL_INST_A2F_R_17_3 (.IN_IBUF(tcdm_rdata_p2[3]),.OUT_IBUF(tcdm_rdata_p2_int[3]));

	IBUF QL_INST_A2F_R_17_4 (.IN_IBUF(tcdm_valid_p2),.OUT_IBUF(tcdm_valid_p2_int));

	IBUF QL_INST_A2F_R_17_5 (.IN_IBUF(tcdm_gnt_p2),.OUT_IBUF(tcdm_gnt_p2_int));

	OBUF QL_INST_F2A_R_18_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[0]),.OUT_OBUF(tcdm_wdata_p2[0]));

	OBUF QL_INST_F2A_R_18_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[1]),.OUT_OBUF(tcdm_wdata_p2[1]));

	OBUF QL_INST_F2A_R_18_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[2]),.OUT_OBUF(tcdm_wdata_p2[2]));

	OBUF QL_INST_F2A_R_18_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[3]),.OUT_OBUF(tcdm_wdata_p2[3]));

	OBUF QL_INST_F2A_R_18_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[4]),.OUT_OBUF(tcdm_wdata_p2[4]));

	OBUF QL_INST_F2A_R_18_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[5]),.OUT_OBUF(tcdm_wdata_p2[5]));

	OBUF QL_INST_F2A_R_18_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[6]),.OUT_OBUF(tcdm_wdata_p2[6]));

	OBUF QL_INST_F2A_R_18_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[7]),.OUT_OBUF(tcdm_wdata_p2[7]));

	OBUF QL_INST_F2A_R_18_9 (.IN_OBUF(tcdm_addr_p2_dup_0[4]),.OUT_OBUF(tcdm_addr_p2[4]));

	OBUF QL_INST_F2A_R_18_10 (.IN_OBUF(tcdm_addr_p2_dup_0[5]),.OUT_OBUF(tcdm_addr_p2[5]));

	OBUF QL_INST_F2A_R_18_11 (.IN_OBUF(tcdm_addr_p2_dup_0[6]),.OUT_OBUF(tcdm_addr_p2[6]));

	OBUF QL_INST_F2A_R_18_12 (.IN_OBUF(tcdm_addr_p2_dup_0[7]),.OUT_OBUF(tcdm_addr_p2[7]));

	OBUF QL_INST_F2A_R_18_13 (.IN_OBUF(tcdm_addr_p2_dup_0[8]),.OUT_OBUF(tcdm_addr_p2[8]));

	OBUF QL_INST_F2A_R_18_14 (.IN_OBUF(tcdm_addr_p2_dup_0[9]),.OUT_OBUF(tcdm_addr_p2[9]));

	IBUF QL_INST_A2F_R_18_0 (.IN_IBUF(tcdm_rdata_p2[4]),.OUT_IBUF(tcdm_rdata_p2_int[4]));

	IBUF QL_INST_A2F_R_18_1 (.IN_IBUF(tcdm_rdata_p2[5]),.OUT_IBUF(tcdm_rdata_p2_int[5]));

	IBUF QL_INST_A2F_R_18_2 (.IN_IBUF(tcdm_rdata_p2[6]),.OUT_IBUF(tcdm_rdata_p2_int[6]));

	IBUF QL_INST_A2F_R_18_3 (.IN_IBUF(tcdm_rdata_p2[7]),.OUT_IBUF(tcdm_rdata_p2_int[7]));

	IBUF QL_INST_A2F_R_18_4 (.IN_IBUF(tcdm_rdata_p2[8]),.OUT_IBUF(tcdm_rdata_p2_int[8]));

	IBUF QL_INST_A2F_R_18_5 (.IN_IBUF(tcdm_rdata_p2[9]),.OUT_IBUF(tcdm_rdata_p2_int[9]));

	IBUF QL_INST_A2F_R_18_6 (.IN_IBUF(tcdm_rdata_p2[10]),.OUT_IBUF(tcdm_rdata_p2_int[10]));

	IBUF QL_INST_A2F_R_18_7 (.IN_IBUF(tcdm_rdata_p2[11]),.OUT_IBUF(tcdm_rdata_p2_int[11]));

	OBUF QL_INST_F2A_R_19_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[8]),.OUT_OBUF(tcdm_wdata_p2[8]));

	OBUF QL_INST_F2A_R_19_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[9]),.OUT_OBUF(tcdm_wdata_p2[9]));

	OBUF QL_INST_F2A_R_19_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[10]),.OUT_OBUF(tcdm_wdata_p2[10]));

	OBUF QL_INST_F2A_R_19_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[11]),.OUT_OBUF(tcdm_wdata_p2[11]));

	OBUF QL_INST_F2A_R_19_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[12]),.OUT_OBUF(tcdm_wdata_p2[12]));

	OBUF QL_INST_F2A_R_19_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[13]),.OUT_OBUF(tcdm_wdata_p2[13]));

	OBUF QL_INST_F2A_R_19_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[14]),.OUT_OBUF(tcdm_wdata_p2[14]));

	OBUF QL_INST_F2A_R_19_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[15]),.OUT_OBUF(tcdm_wdata_p2[15]));

	OBUF QL_INST_F2A_R_19_8 (.IN_OBUF(tcdm_addr_p2_dup_0[10]),.OUT_OBUF(tcdm_addr_p2[10]));

	OBUF QL_INST_F2A_R_19_9 (.IN_OBUF(tcdm_addr_p2_dup_0[11]),.OUT_OBUF(tcdm_addr_p2[11]));

	OBUF QL_INST_F2A_R_19_10 (.IN_OBUF(tcdm_addr_p2_dup_0[12]),.OUT_OBUF(tcdm_addr_p2[12]));

	OBUF QL_INST_F2A_R_19_11 (.IN_OBUF(tcdm_addr_p2_dup_0[13]),.OUT_OBUF(tcdm_addr_p2[13]));

	IBUF QL_INST_A2F_R_19_0 (.IN_IBUF(tcdm_rdata_p2[12]),.OUT_IBUF(tcdm_rdata_p2_int[12]));

	IBUF QL_INST_A2F_R_19_1 (.IN_IBUF(tcdm_rdata_p2[13]),.OUT_IBUF(tcdm_rdata_p2_int[13]));

	IBUF QL_INST_A2F_R_19_2 (.IN_IBUF(tcdm_rdata_p2[14]),.OUT_IBUF(tcdm_rdata_p2_int[14]));

	IBUF QL_INST_A2F_R_19_3 (.IN_IBUF(tcdm_rdata_p2[15]),.OUT_IBUF(tcdm_rdata_p2_int[15]));

	OBUF QL_INST_F2A_R_20_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[16]),.OUT_OBUF(tcdm_wdata_p2[16]));

	OBUF QL_INST_F2A_R_20_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[17]),.OUT_OBUF(tcdm_wdata_p2[17]));

	OBUF QL_INST_F2A_R_20_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[18]),.OUT_OBUF(tcdm_wdata_p2[18]));

	OBUF QL_INST_F2A_R_20_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[19]),.OUT_OBUF(tcdm_wdata_p2[19]));

	OBUF QL_INST_F2A_R_20_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[20]),.OUT_OBUF(tcdm_wdata_p2[20]));

	OBUF QL_INST_F2A_R_20_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[21]),.OUT_OBUF(tcdm_wdata_p2[21]));

	OBUF QL_INST_F2A_R_20_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[22]),.OUT_OBUF(tcdm_wdata_p2[22]));

	OBUF QL_INST_F2A_R_20_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[23]),.OUT_OBUF(tcdm_wdata_p2[23]));

	OBUF QL_INST_F2A_R_20_12 (.IN_OBUF(tcdm_addr_p2_dup_0[14]),.OUT_OBUF(tcdm_addr_p2[14]));

	OBUF QL_INST_F2A_R_20_13 (.IN_OBUF(tcdm_addr_p2_dup_0[15]),.OUT_OBUF(tcdm_addr_p2[15]));

	OBUF QL_INST_F2A_R_20_14 (.IN_OBUF(tcdm_addr_p2_dup_0[16]),.OUT_OBUF(tcdm_addr_p2[16]));

	OBUF QL_INST_F2A_R_20_15 (.IN_OBUF(tcdm_addr_p2_dup_0[17]),.OUT_OBUF(tcdm_addr_p2[17]));

	OBUF QL_INST_F2A_R_20_16 (.IN_OBUF(tcdm_addr_p2_dup_0[18]),.OUT_OBUF(tcdm_addr_p2[18]));

	OBUF QL_INST_F2A_R_20_17 (.IN_OBUF(tcdm_addr_p2_dup_0[19]),.OUT_OBUF(tcdm_addr_p2[19]));

	IBUF QL_INST_A2F_R_20_1 (.IN_IBUF(tcdm_rdata_p2[16]),.OUT_IBUF(tcdm_rdata_p2_int[16]));

	IBUF QL_INST_A2F_R_20_2 (.IN_IBUF(tcdm_rdata_p2[17]),.OUT_IBUF(tcdm_rdata_p2_int[17]));

	IBUF QL_INST_A2F_R_20_3 (.IN_IBUF(tcdm_rdata_p2[18]),.OUT_IBUF(tcdm_rdata_p2_int[18]));

	IBUF QL_INST_A2F_R_20_4 (.IN_IBUF(tcdm_rdata_p2[19]),.OUT_IBUF(tcdm_rdata_p2_int[19]));

	IBUF QL_INST_A2F_R_20_5 (.IN_IBUF(tcdm_rdata_p2[20]),.OUT_IBUF(tcdm_rdata_p2_int[20]));

	IBUF QL_INST_A2F_R_20_6 (.IN_IBUF(tcdm_rdata_p2[21]),.OUT_IBUF(tcdm_rdata_p2_int[21]));

	OBUF QL_INST_F2A_R_21_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[24]),.OUT_OBUF(tcdm_wdata_p2[24]));

	OBUF QL_INST_F2A_R_21_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[25]),.OUT_OBUF(tcdm_wdata_p2[25]));

	OBUF QL_INST_F2A_R_21_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[26]),.OUT_OBUF(tcdm_wdata_p2[26]));

	OBUF QL_INST_F2A_R_21_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[27]),.OUT_OBUF(tcdm_wdata_p2[27]));

	OBUF QL_INST_F2A_R_21_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[28]),.OUT_OBUF(tcdm_wdata_p2[28]));

	OBUF QL_INST_F2A_R_21_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[29]),.OUT_OBUF(tcdm_wdata_p2[29]));

	OBUF QL_INST_F2A_R_21_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[30]),.OUT_OBUF(tcdm_wdata_p2[30]));

	OBUF QL_INST_F2A_R_21_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[31]),.OUT_OBUF(tcdm_wdata_p2[31]));

	IBUF QL_INST_A2F_R_21_0 (.IN_IBUF(tcdm_rdata_p2[22]),.OUT_IBUF(tcdm_rdata_p2_int[22]));

	IBUF QL_INST_A2F_R_21_1 (.IN_IBUF(tcdm_rdata_p2[23]),.OUT_IBUF(tcdm_rdata_p2_int[23]));

	IBUF QL_INST_A2F_R_21_2 (.IN_IBUF(tcdm_rdata_p2[24]),.OUT_IBUF(tcdm_rdata_p2_int[24]));

	IBUF QL_INST_A2F_R_21_3 (.IN_IBUF(tcdm_rdata_p2[25]),.OUT_IBUF(tcdm_rdata_p2_int[25]));

	IBUF QL_INST_A2F_R_21_4 (.IN_IBUF(tcdm_rdata_p2[26]),.OUT_IBUF(tcdm_rdata_p2_int[26]));

	IBUF QL_INST_A2F_R_21_5 (.IN_IBUF(tcdm_rdata_p2[27]),.OUT_IBUF(tcdm_rdata_p2_int[27]));

	IBUF QL_INST_A2F_R_22_0 (.IN_IBUF(tcdm_rdata_p2[28]),.OUT_IBUF(tcdm_rdata_p2_int[28]));

	IBUF QL_INST_A2F_R_22_1 (.IN_IBUF(tcdm_rdata_p2[29]),.OUT_IBUF(tcdm_rdata_p2_int[29]));

	IBUF QL_INST_A2F_R_22_2 (.IN_IBUF(tcdm_rdata_p2[30]),.OUT_IBUF(tcdm_rdata_p2_int[30]));

	IBUF QL_INST_A2F_R_22_3 (.IN_IBUF(tcdm_rdata_p2[31]),.OUT_IBUF(tcdm_rdata_p2_int[31]));

	OBUF QL_INST_F2A_R_23_0 (.IN_OBUF(CLK_int_0__CAND0_BRSTR_33_padClk),.OUT_OBUF(tcdm_clk_p3));

	OBUF QL_INST_F2A_R_23_1 (.IN_OBUF(tcdm_req_p3_dup_0),.OUT_OBUF(tcdm_req_p3));

	OBUF QL_INST_F2A_R_23_2 (.IN_OBUF(tcdm_wen_p3_dup_0),.OUT_OBUF(tcdm_wen_p3));

	OBUF QL_INST_F2A_R_23_3 (.IN_OBUF(tcdm_be_p3_dup_0[0]),.OUT_OBUF(tcdm_be_p3[0]));

	OBUF QL_INST_F2A_R_23_4 (.IN_OBUF(tcdm_be_p3_dup_0[1]),.OUT_OBUF(tcdm_be_p3[1]));

	OBUF QL_INST_F2A_R_23_5 (.IN_OBUF(tcdm_be_p3_dup_0[2]),.OUT_OBUF(tcdm_be_p3[2]));

	OBUF QL_INST_F2A_R_23_6 (.IN_OBUF(tcdm_be_p3_dup_0[3]),.OUT_OBUF(tcdm_be_p3[3]));

	OBUF QL_INST_F2A_R_23_8 (.IN_OBUF(tcdm_addr_p3_dup_0[0]),.OUT_OBUF(tcdm_addr_p3[0]));

	OBUF QL_INST_F2A_R_23_9 (.IN_OBUF(tcdm_addr_p3_dup_0[1]),.OUT_OBUF(tcdm_addr_p3[1]));

	OBUF QL_INST_F2A_R_23_10 (.IN_OBUF(tcdm_addr_p3_dup_0[2]),.OUT_OBUF(tcdm_addr_p3[2]));

	OBUF QL_INST_F2A_R_23_11 (.IN_OBUF(tcdm_addr_p3_dup_0[3]),.OUT_OBUF(tcdm_addr_p3[3]));

	IBUF QL_INST_A2F_R_23_0 (.IN_IBUF(tcdm_rdata_p3[0]),.OUT_IBUF(tcdm_rdata_p3_int[0]));

	IBUF QL_INST_A2F_R_23_1 (.IN_IBUF(tcdm_rdata_p3[1]),.OUT_IBUF(tcdm_rdata_p3_int[1]));

	IBUF QL_INST_A2F_R_23_2 (.IN_IBUF(tcdm_rdata_p3[2]),.OUT_IBUF(tcdm_rdata_p3_int[2]));

	IBUF QL_INST_A2F_R_23_3 (.IN_IBUF(tcdm_rdata_p3[3]),.OUT_IBUF(tcdm_rdata_p3_int[3]));

	IBUF QL_INST_A2F_R_23_4 (.IN_IBUF(tcdm_valid_p3),.OUT_IBUF(tcdm_valid_p3_int));

	IBUF QL_INST_A2F_R_23_5 (.IN_IBUF(tcdm_gnt_p3),.OUT_IBUF(tcdm_gnt_p3_int));

	OBUF QL_INST_F2A_R_24_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[0]),.OUT_OBUF(tcdm_wdata_p3[0]));

	OBUF QL_INST_F2A_R_24_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[1]),.OUT_OBUF(tcdm_wdata_p3[1]));

	OBUF QL_INST_F2A_R_24_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[2]),.OUT_OBUF(tcdm_wdata_p3[2]));

	OBUF QL_INST_F2A_R_24_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[3]),.OUT_OBUF(tcdm_wdata_p3[3]));

	OBUF QL_INST_F2A_R_24_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[4]),.OUT_OBUF(tcdm_wdata_p3[4]));

	OBUF QL_INST_F2A_R_24_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[5]),.OUT_OBUF(tcdm_wdata_p3[5]));

	OBUF QL_INST_F2A_R_24_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[6]),.OUT_OBUF(tcdm_wdata_p3[6]));

	OBUF QL_INST_F2A_R_24_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[7]),.OUT_OBUF(tcdm_wdata_p3[7]));

	OBUF QL_INST_F2A_R_24_9 (.IN_OBUF(tcdm_addr_p3_dup_0[4]),.OUT_OBUF(tcdm_addr_p3[4]));

	OBUF QL_INST_F2A_R_24_10 (.IN_OBUF(tcdm_addr_p3_dup_0[5]),.OUT_OBUF(tcdm_addr_p3[5]));

	OBUF QL_INST_F2A_R_24_11 (.IN_OBUF(tcdm_addr_p3_dup_0[6]),.OUT_OBUF(tcdm_addr_p3[6]));

	OBUF QL_INST_F2A_R_24_12 (.IN_OBUF(tcdm_addr_p3_dup_0[7]),.OUT_OBUF(tcdm_addr_p3[7]));

	OBUF QL_INST_F2A_R_24_13 (.IN_OBUF(tcdm_addr_p3_dup_0[8]),.OUT_OBUF(tcdm_addr_p3[8]));

	OBUF QL_INST_F2A_R_24_14 (.IN_OBUF(tcdm_addr_p3_dup_0[9]),.OUT_OBUF(tcdm_addr_p3[9]));

	IBUF QL_INST_A2F_R_24_0 (.IN_IBUF(tcdm_rdata_p3[4]),.OUT_IBUF(tcdm_rdata_p3_int[4]));

	IBUF QL_INST_A2F_R_24_1 (.IN_IBUF(tcdm_rdata_p3[5]),.OUT_IBUF(tcdm_rdata_p3_int[5]));

	IBUF QL_INST_A2F_R_24_2 (.IN_IBUF(tcdm_rdata_p3[6]),.OUT_IBUF(tcdm_rdata_p3_int[6]));

	IBUF QL_INST_A2F_R_24_3 (.IN_IBUF(tcdm_rdata_p3[7]),.OUT_IBUF(tcdm_rdata_p3_int[7]));

	IBUF QL_INST_A2F_R_24_4 (.IN_IBUF(tcdm_rdata_p3[8]),.OUT_IBUF(tcdm_rdata_p3_int[8]));

	IBUF QL_INST_A2F_R_24_5 (.IN_IBUF(tcdm_rdata_p3[9]),.OUT_IBUF(tcdm_rdata_p3_int[9]));

	IBUF QL_INST_A2F_R_24_6 (.IN_IBUF(tcdm_rdata_p3[10]),.OUT_IBUF(tcdm_rdata_p3_int[10]));

	IBUF QL_INST_A2F_R_24_7 (.IN_IBUF(tcdm_rdata_p3[11]),.OUT_IBUF(tcdm_rdata_p3_int[11]));

	OBUF QL_INST_F2A_R_25_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[8]),.OUT_OBUF(tcdm_wdata_p3[8]));

	OBUF QL_INST_F2A_R_25_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[9]),.OUT_OBUF(tcdm_wdata_p3[9]));

	OBUF QL_INST_F2A_R_25_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[10]),.OUT_OBUF(tcdm_wdata_p3[10]));

	OBUF QL_INST_F2A_R_25_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[11]),.OUT_OBUF(tcdm_wdata_p3[11]));

	OBUF QL_INST_F2A_R_25_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[12]),.OUT_OBUF(tcdm_wdata_p3[12]));

	OBUF QL_INST_F2A_R_25_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[13]),.OUT_OBUF(tcdm_wdata_p3[13]));

	OBUF QL_INST_F2A_R_25_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[14]),.OUT_OBUF(tcdm_wdata_p3[14]));

	OBUF QL_INST_F2A_R_25_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[15]),.OUT_OBUF(tcdm_wdata_p3[15]));

	OBUF QL_INST_F2A_R_25_8 (.IN_OBUF(tcdm_addr_p3_dup_0[10]),.OUT_OBUF(tcdm_addr_p3[10]));

	OBUF QL_INST_F2A_R_25_9 (.IN_OBUF(tcdm_addr_p3_dup_0[11]),.OUT_OBUF(tcdm_addr_p3[11]));

	OBUF QL_INST_F2A_R_25_10 (.IN_OBUF(tcdm_addr_p3_dup_0[12]),.OUT_OBUF(tcdm_addr_p3[12]));

	OBUF QL_INST_F2A_R_25_11 (.IN_OBUF(tcdm_addr_p3_dup_0[13]),.OUT_OBUF(tcdm_addr_p3[13]));

	IBUF QL_INST_A2F_R_25_0 (.IN_IBUF(tcdm_rdata_p3[12]),.OUT_IBUF(tcdm_rdata_p3_int[12]));

	IBUF QL_INST_A2F_R_25_1 (.IN_IBUF(tcdm_rdata_p3[13]),.OUT_IBUF(tcdm_rdata_p3_int[13]));

	IBUF QL_INST_A2F_R_25_2 (.IN_IBUF(tcdm_rdata_p3[14]),.OUT_IBUF(tcdm_rdata_p3_int[14]));

	IBUF QL_INST_A2F_R_25_3 (.IN_IBUF(tcdm_rdata_p3[15]),.OUT_IBUF(tcdm_rdata_p3_int[15]));

	OBUF QL_INST_F2A_R_26_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[16]),.OUT_OBUF(tcdm_wdata_p3[16]));

	OBUF QL_INST_F2A_R_26_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[17]),.OUT_OBUF(tcdm_wdata_p3[17]));

	OBUF QL_INST_F2A_R_26_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[18]),.OUT_OBUF(tcdm_wdata_p3[18]));

	OBUF QL_INST_F2A_R_26_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[19]),.OUT_OBUF(tcdm_wdata_p3[19]));

	OBUF QL_INST_F2A_R_26_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[20]),.OUT_OBUF(tcdm_wdata_p3[20]));

	OBUF QL_INST_F2A_R_26_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[21]),.OUT_OBUF(tcdm_wdata_p3[21]));

	OBUF QL_INST_F2A_R_26_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[22]),.OUT_OBUF(tcdm_wdata_p3[22]));

	OBUF QL_INST_F2A_R_26_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[23]),.OUT_OBUF(tcdm_wdata_p3[23]));

	OBUF QL_INST_F2A_R_26_12 (.IN_OBUF(tcdm_addr_p3_dup_0[14]),.OUT_OBUF(tcdm_addr_p3[14]));

	OBUF QL_INST_F2A_R_26_13 (.IN_OBUF(tcdm_addr_p3_dup_0[15]),.OUT_OBUF(tcdm_addr_p3[15]));

	OBUF QL_INST_F2A_R_26_14 (.IN_OBUF(tcdm_addr_p3_dup_0[16]),.OUT_OBUF(tcdm_addr_p3[16]));

	OBUF QL_INST_F2A_R_26_15 (.IN_OBUF(tcdm_addr_p3_dup_0[17]),.OUT_OBUF(tcdm_addr_p3[17]));

	OBUF QL_INST_F2A_R_26_16 (.IN_OBUF(tcdm_addr_p3_dup_0[18]),.OUT_OBUF(tcdm_addr_p3[18]));

	OBUF QL_INST_F2A_R_26_17 (.IN_OBUF(tcdm_addr_p3_dup_0[19]),.OUT_OBUF(tcdm_addr_p3[19]));

	IBUF QL_INST_A2F_R_26_1 (.IN_IBUF(tcdm_rdata_p3[16]),.OUT_IBUF(tcdm_rdata_p3_int[16]));

	IBUF QL_INST_A2F_R_26_2 (.IN_IBUF(tcdm_rdata_p3[17]),.OUT_IBUF(tcdm_rdata_p3_int[17]));

	IBUF QL_INST_A2F_R_26_3 (.IN_IBUF(tcdm_rdata_p3[18]),.OUT_IBUF(tcdm_rdata_p3_int[18]));

	IBUF QL_INST_A2F_R_26_4 (.IN_IBUF(tcdm_rdata_p3[19]),.OUT_IBUF(tcdm_rdata_p3_int[19]));

	IBUF QL_INST_A2F_R_26_5 (.IN_IBUF(tcdm_rdata_p3[20]),.OUT_IBUF(tcdm_rdata_p3_int[20]));

	IBUF QL_INST_A2F_R_26_6 (.IN_IBUF(tcdm_rdata_p3[21]),.OUT_IBUF(tcdm_rdata_p3_int[21]));

	OBUF QL_INST_F2A_R_27_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[24]),.OUT_OBUF(tcdm_wdata_p3[24]));

	OBUF QL_INST_F2A_R_27_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[25]),.OUT_OBUF(tcdm_wdata_p3[25]));

	OBUF QL_INST_F2A_R_27_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[26]),.OUT_OBUF(tcdm_wdata_p3[26]));

	OBUF QL_INST_F2A_R_27_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[27]),.OUT_OBUF(tcdm_wdata_p3[27]));

	OBUF QL_INST_F2A_R_27_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[28]),.OUT_OBUF(tcdm_wdata_p3[28]));

	OBUF QL_INST_F2A_R_27_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[29]),.OUT_OBUF(tcdm_wdata_p3[29]));

	OBUF QL_INST_F2A_R_27_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[30]),.OUT_OBUF(tcdm_wdata_p3[30]));

	OBUF QL_INST_F2A_R_27_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[31]),.OUT_OBUF(tcdm_wdata_p3[31]));

	IBUF QL_INST_A2F_R_27_0 (.IN_IBUF(tcdm_rdata_p3[22]),.OUT_IBUF(tcdm_rdata_p3_int[22]));

	IBUF QL_INST_A2F_R_27_1 (.IN_IBUF(tcdm_rdata_p3[23]),.OUT_IBUF(tcdm_rdata_p3_int[23]));

	IBUF QL_INST_A2F_R_27_2 (.IN_IBUF(tcdm_rdata_p3[24]),.OUT_IBUF(tcdm_rdata_p3_int[24]));

	IBUF QL_INST_A2F_R_27_3 (.IN_IBUF(tcdm_rdata_p3[25]),.OUT_IBUF(tcdm_rdata_p3_int[25]));

	IBUF QL_INST_A2F_R_27_4 (.IN_IBUF(tcdm_rdata_p3[26]),.OUT_IBUF(tcdm_rdata_p3_int[26]));

	IBUF QL_INST_A2F_R_27_5 (.IN_IBUF(tcdm_rdata_p3[27]),.OUT_IBUF(tcdm_rdata_p3_int[27]));

	IBUF QL_INST_A2F_R_28_0 (.IN_IBUF(tcdm_rdata_p3[28]),.OUT_IBUF(tcdm_rdata_p3_int[28]));

	IBUF QL_INST_A2F_R_28_1 (.IN_IBUF(tcdm_rdata_p3[29]),.OUT_IBUF(tcdm_rdata_p3_int[29]));

	IBUF QL_INST_A2F_R_28_2 (.IN_IBUF(tcdm_rdata_p3[30]),.OUT_IBUF(tcdm_rdata_p3_int[30]));

	IBUF QL_INST_A2F_R_28_3 (.IN_IBUF(tcdm_rdata_p3[31]),.OUT_IBUF(tcdm_rdata_p3_int[31]));

	IBUF QL_INST_A2F_R_29_2 (.IN_IBUF(RESET[1]),.OUT_IBUF(RESET_int[1]));

	OBUF QL_INST_F2A_B_2_0 (.IN_OBUF(CLK_int_0__CAND0_BLSBL_2_padClk),.OUT_OBUF(m1_oper0_wclk));

	OBUF QL_INST_F2A_B_2_1 (.IN_OBUF(m0_oper0_wmode_dup_0[1]),.OUT_OBUF(m1_oper0_wmode[1]));

	OBUF QL_INST_F2A_B_2_2 (.IN_OBUF(m0_oper0_wmode_dup_0[0]),.OUT_OBUF(m1_oper0_wmode[0]));

	OBUF QL_INST_F2A_B_2_3 (.IN_OBUF(m0_oper0_wdsel_dup_0),.OUT_OBUF(m1_oper0_wdsel));

	OBUF QL_INST_F2A_B_2_4 (.IN_OBUF(m0_oper0_rmode_dup_0[1]),.OUT_OBUF(m1_oper0_rmode[1]));

	OBUF QL_INST_F2A_B_2_5 (.IN_OBUF(m0_oper0_rmode_dup_0[0]),.OUT_OBUF(m1_oper0_rmode[0]));

	OBUF QL_INST_F2A_B_2_6 (.IN_OBUF(m1_oper0_wdata_dup_0[31]),.OUT_OBUF(m1_oper0_wdata[31]));

	OBUF QL_INST_F2A_B_2_7 (.IN_OBUF(m1_oper0_wdata_dup_0[30]),.OUT_OBUF(m1_oper0_wdata[30]));

	OBUF QL_INST_F2A_B_2_8 (.IN_OBUF(m1_oper0_wdata_dup_0[29]),.OUT_OBUF(m1_oper0_wdata[29]));

	OBUF QL_INST_F2A_B_2_9 (.IN_OBUF(m1_oper0_wdata_dup_0[28]),.OUT_OBUF(m1_oper0_wdata[28]));

	OBUF QL_INST_F2A_B_2_10 (.IN_OBUF(m1_oper0_wdata_dup_0[27]),.OUT_OBUF(m1_oper0_wdata[27]));

	OBUF QL_INST_F2A_B_2_11 (.IN_OBUF(m1_oper0_wdata_dup_0[26]),.OUT_OBUF(m1_oper0_wdata[26]));

	OBUF QL_INST_F2A_B_2_12 (.IN_OBUF(m1_oper0_wdata_dup_0[25]),.OUT_OBUF(m1_oper0_wdata[25]));

	OBUF QL_INST_F2A_B_2_13 (.IN_OBUF(m1_oper0_wdata_dup_0[24]),.OUT_OBUF(m1_oper0_wdata[24]));

	OBUF QL_INST_F2A_B_2_14 (.IN_OBUF(m1_oper0_wdata_dup_0[23]),.OUT_OBUF(m1_oper0_wdata[23]));

	OBUF QL_INST_F2A_B_2_15 (.IN_OBUF(m1_oper0_wdata_dup_0[22]),.OUT_OBUF(m1_oper0_wdata[22]));

	OBUF QL_INST_F2A_B_2_16 (.IN_OBUF(m1_oper0_wdata_dup_0[21]),.OUT_OBUF(m1_oper0_wdata[21]));

	OBUF QL_INST_F2A_B_2_17 (.IN_OBUF(m1_oper0_wdata_dup_0[20]),.OUT_OBUF(m1_oper0_wdata[20]));

	IBUF QL_INST_A2F_B_2_0 (.IN_IBUF(m1_oper0_rdata[31]),.OUT_IBUF(m1_oper0_rdata_int[31]));

	IBUF QL_INST_A2F_B_2_1 (.IN_IBUF(m1_oper0_rdata[30]),.OUT_IBUF(m1_oper0_rdata_int[30]));

	IBUF QL_INST_A2F_B_2_2 (.IN_IBUF(m1_oper0_rdata[29]),.OUT_IBUF(m1_oper0_rdata_int[29]));

	IBUF QL_INST_A2F_B_2_3 (.IN_IBUF(m1_oper0_rdata[28]),.OUT_IBUF(m1_oper0_rdata_int[28]));

	OBUF QL_INST_F2A_B_3_0 (.IN_OBUF(m1_oper0_wdata_dup_0[19]),.OUT_OBUF(m1_oper0_wdata[19]));

	OBUF QL_INST_F2A_B_3_1 (.IN_OBUF(m1_oper0_wdata_dup_0[18]),.OUT_OBUF(m1_oper0_wdata[18]));

	OBUF QL_INST_F2A_B_3_2 (.IN_OBUF(m1_oper0_wdata_dup_0[17]),.OUT_OBUF(m1_oper0_wdata[17]));

	OBUF QL_INST_F2A_B_3_3 (.IN_OBUF(m1_oper0_wdata_dup_0[16]),.OUT_OBUF(m1_oper0_wdata[16]));

	OBUF QL_INST_F2A_B_3_4 (.IN_OBUF(m1_oper0_wdata_dup_0[15]),.OUT_OBUF(m1_oper0_wdata[15]));

	OBUF QL_INST_F2A_B_3_5 (.IN_OBUF(m1_oper0_wdata_dup_0[14]),.OUT_OBUF(m1_oper0_wdata[14]));

	OBUF QL_INST_F2A_B_3_6 (.IN_OBUF(m1_oper0_wdata_dup_0[13]),.OUT_OBUF(m1_oper0_wdata[13]));

	OBUF QL_INST_F2A_B_3_7 (.IN_OBUF(m1_oper0_wdata_dup_0[12]),.OUT_OBUF(m1_oper0_wdata[12]));

	OBUF QL_INST_F2A_B_3_8 (.IN_OBUF(m1_oper0_wdata_dup_0[11]),.OUT_OBUF(m1_oper0_wdata[11]));

	OBUF QL_INST_F2A_B_3_9 (.IN_OBUF(m1_oper0_wdata_dup_0[10]),.OUT_OBUF(m1_oper0_wdata[10]));

	OBUF QL_INST_F2A_B_3_10 (.IN_OBUF(m1_oper0_wdata_dup_0[9]),.OUT_OBUF(m1_oper0_wdata[9]));

	OBUF QL_INST_F2A_B_3_11 (.IN_OBUF(m1_oper0_wdata_dup_0[8]),.OUT_OBUF(m1_oper0_wdata[8]));

	IBUF QL_INST_A2F_B_3_0 (.IN_IBUF(m1_oper0_rdata[27]),.OUT_IBUF(m1_oper0_rdata_int[27]));

	IBUF QL_INST_A2F_B_3_1 (.IN_IBUF(m1_oper0_rdata[26]),.OUT_IBUF(m1_oper0_rdata_int[26]));

	IBUF QL_INST_A2F_B_3_2 (.IN_IBUF(m1_oper0_rdata[25]),.OUT_IBUF(m1_oper0_rdata_int[25]));

	IBUF QL_INST_A2F_B_3_3 (.IN_IBUF(m1_oper0_rdata[24]),.OUT_IBUF(m1_oper0_rdata_int[24]));

	IBUF QL_INST_A2F_B_3_4 (.IN_IBUF(m1_oper0_rdata[23]),.OUT_IBUF(m1_oper0_rdata_int[23]));

	IBUF QL_INST_A2F_B_3_5 (.IN_IBUF(m1_oper0_rdata[22]),.OUT_IBUF(m1_oper0_rdata_int[22]));

	OBUF QL_INST_F2A_B_4_0 (.IN_OBUF(m1_oper0_wdata_dup_0[7]),.OUT_OBUF(m1_oper0_wdata[7]));

	OBUF QL_INST_F2A_B_4_1 (.IN_OBUF(m1_oper0_wdata_dup_0[6]),.OUT_OBUF(m1_oper0_wdata[6]));

	OBUF QL_INST_F2A_B_4_2 (.IN_OBUF(m1_oper0_wdata_dup_0[5]),.OUT_OBUF(m1_oper0_wdata[5]));

	OBUF QL_INST_F2A_B_4_3 (.IN_OBUF(m1_oper0_wdata_dup_0[4]),.OUT_OBUF(m1_oper0_wdata[4]));

	OBUF QL_INST_F2A_B_4_4 (.IN_OBUF(m1_oper0_wdata_dup_0[3]),.OUT_OBUF(m1_oper0_wdata[3]));

	OBUF QL_INST_F2A_B_4_5 (.IN_OBUF(m1_oper0_wdata_dup_0[2]),.OUT_OBUF(m1_oper0_wdata[2]));

	OBUF QL_INST_F2A_B_4_6 (.IN_OBUF(m1_oper0_wdata_dup_0[1]),.OUT_OBUF(m1_oper0_wdata[1]));

	OBUF QL_INST_F2A_B_4_7 (.IN_OBUF(m1_oper0_wdata_dup_0[0]),.OUT_OBUF(m1_oper0_wdata[0]));

	OBUF QL_INST_F2A_B_4_8 (.IN_OBUF(m1_oper0_waddr_dup_0[11]),.OUT_OBUF(m1_oper0_waddr[11]));

	OBUF QL_INST_F2A_B_4_9 (.IN_OBUF(m1_oper0_waddr_dup_0[10]),.OUT_OBUF(m1_oper0_waddr[10]));

	OBUF QL_INST_F2A_B_4_10 (.IN_OBUF(m1_oper0_waddr_dup_0[9]),.OUT_OBUF(m1_oper0_waddr[9]));

	OBUF QL_INST_F2A_B_4_11 (.IN_OBUF(m1_oper0_waddr_dup_0[8]),.OUT_OBUF(m1_oper0_waddr[8]));

	OBUF QL_INST_F2A_B_4_12 (.IN_OBUF(m1_oper0_waddr_dup_0[7]),.OUT_OBUF(m1_oper0_waddr[7]));

	OBUF QL_INST_F2A_B_4_13 (.IN_OBUF(m1_oper0_waddr_dup_0[6]),.OUT_OBUF(m1_oper0_waddr[6]));

	OBUF QL_INST_F2A_B_4_14 (.IN_OBUF(m1_oper0_waddr_dup_0[5]),.OUT_OBUF(m1_oper0_waddr[5]));

	OBUF QL_INST_F2A_B_4_15 (.IN_OBUF(m1_oper0_waddr_dup_0[4]),.OUT_OBUF(m1_oper0_waddr[4]));

	OBUF QL_INST_F2A_B_4_16 (.IN_OBUF(m1_oper0_waddr_dup_0[3]),.OUT_OBUF(m1_oper0_waddr[3]));

	OBUF QL_INST_F2A_B_4_17 (.IN_OBUF(m1_oper0_waddr_dup_0[2]),.OUT_OBUF(m1_oper0_waddr[2]));

	IBUF QL_INST_A2F_B_4_0 (.IN_IBUF(m1_oper0_rdata[21]),.OUT_IBUF(m1_oper0_rdata_int[21]));

	IBUF QL_INST_A2F_B_4_1 (.IN_IBUF(m1_oper0_rdata[20]),.OUT_IBUF(m1_oper0_rdata_int[20]));

	IBUF QL_INST_A2F_B_4_2 (.IN_IBUF(m1_oper0_rdata[19]),.OUT_IBUF(m1_oper0_rdata_int[19]));

	IBUF QL_INST_A2F_B_4_3 (.IN_IBUF(m1_oper0_rdata[18]),.OUT_IBUF(m1_oper0_rdata_int[18]));

	IBUF QL_INST_A2F_B_4_4 (.IN_IBUF(m1_oper0_rdata[17]),.OUT_IBUF(m1_oper0_rdata_int[17]));

	IBUF QL_INST_A2F_B_4_5 (.IN_IBUF(m1_oper0_rdata[16]),.OUT_IBUF(m1_oper0_rdata_int[16]));

	IBUF QL_INST_A2F_B_4_6 (.IN_IBUF(m1_oper0_rdata[15]),.OUT_IBUF(m1_oper0_rdata_int[15]));

	IBUF QL_INST_A2F_B_4_7 (.IN_IBUF(m1_oper0_rdata[14]),.OUT_IBUF(m1_oper0_rdata_int[14]));

	OBUF QL_INST_F2A_B_5_0 (.IN_OBUF(m1_oper0_waddr_dup_0[1]),.OUT_OBUF(m1_oper0_waddr[1]));

	OBUF QL_INST_F2A_B_5_1 (.IN_OBUF(m1_oper0_waddr_dup_0[0]),.OUT_OBUF(m1_oper0_waddr[0]));

	OBUF QL_INST_F2A_B_5_2 (.IN_OBUF(m1_oper0_we_dup_0),.OUT_OBUF(m1_oper0_we));

	OBUF QL_INST_F2A_B_5_3 (.IN_OBUF(m1_oper0_raddr_dup_0[11]),.OUT_OBUF(m1_oper0_raddr[11]));

	OBUF QL_INST_F2A_B_5_4 (.IN_OBUF(m1_oper0_raddr_dup_0[10]),.OUT_OBUF(m1_oper0_raddr[10]));

	OBUF QL_INST_F2A_B_5_5 (.IN_OBUF(m1_oper0_raddr_dup_0[9]),.OUT_OBUF(m1_oper0_raddr[9]));

	OBUF QL_INST_F2A_B_5_6 (.IN_OBUF(m1_oper0_raddr_dup_0[8]),.OUT_OBUF(m1_oper0_raddr[8]));

	OBUF QL_INST_F2A_B_5_7 (.IN_OBUF(m1_oper0_raddr_dup_0[7]),.OUT_OBUF(m1_oper0_raddr[7]));

	OBUF QL_INST_F2A_B_5_8 (.IN_OBUF(m1_oper0_raddr_dup_0[6]),.OUT_OBUF(m1_oper0_raddr[6]));

	OBUF QL_INST_F2A_B_5_9 (.IN_OBUF(m1_oper0_raddr_dup_0[5]),.OUT_OBUF(m1_oper0_raddr[5]));

	OBUF QL_INST_F2A_B_5_10 (.IN_OBUF(m1_oper0_raddr_dup_0[4]),.OUT_OBUF(m1_oper0_raddr[4]));

	OBUF QL_INST_F2A_B_5_11 (.IN_OBUF(m1_oper0_raddr_dup_0[3]),.OUT_OBUF(m1_oper0_raddr[3]));

	IBUF QL_INST_A2F_B_5_0 (.IN_IBUF(m1_oper0_rdata[13]),.OUT_IBUF(m1_oper0_rdata_int[13]));

	IBUF QL_INST_A2F_B_5_1 (.IN_IBUF(m1_oper0_rdata[12]),.OUT_IBUF(m1_oper0_rdata_int[12]));

	IBUF QL_INST_A2F_B_5_2 (.IN_IBUF(m1_oper0_rdata[11]),.OUT_IBUF(m1_oper0_rdata_int[11]));

	IBUF QL_INST_A2F_B_5_3 (.IN_IBUF(m1_oper0_rdata[10]),.OUT_IBUF(m1_oper0_rdata_int[10]));

	IBUF QL_INST_A2F_B_5_4 (.IN_IBUF(m1_oper0_rdata[9]),.OUT_IBUF(m1_oper0_rdata_int[9]));

	IBUF QL_INST_A2F_B_5_5 (.IN_IBUF(m1_oper0_rdata[8]),.OUT_IBUF(m1_oper0_rdata_int[8]));

	OBUF QL_INST_F2A_B_6_0 (.IN_OBUF(CLK_int_0__CAND0_BLSBL_6_padClk),.OUT_OBUF(m1_oper0_rclk));

	OBUF QL_INST_F2A_B_6_1 (.IN_OBUF(m1_oper0_raddr_dup_0[2]),.OUT_OBUF(m1_oper0_raddr[2]));

	OBUF QL_INST_F2A_B_6_2 (.IN_OBUF(m1_oper0_raddr_dup_0[1]),.OUT_OBUF(m1_oper0_raddr[1]));

	OBUF QL_INST_F2A_B_6_3 (.IN_OBUF(m1_oper0_raddr_dup_0[0]),.OUT_OBUF(m1_oper0_raddr[0]));

	OBUF QL_INST_F2A_B_6_4 (.IN_OBUF(m1_m0_osel_dup_0),.OUT_OBUF(m1_m0_osel));

	OBUF QL_INST_F2A_B_6_5 (.IN_OBUF(m1_m0_clken_dup_0),.OUT_OBUF(m1_m0_clken));

	OBUF QL_INST_F2A_B_6_6 (.IN_OBUF(m1_m0_outsel_dup_0[5]),.OUT_OBUF(m1_m0_outsel[5]));

	OBUF QL_INST_F2A_B_6_7 (.IN_OBUF(m1_m0_outsel_dup_0[4]),.OUT_OBUF(m1_m0_outsel[4]));

	OBUF QL_INST_F2A_B_6_8 (.IN_OBUF(m1_m0_outsel_dup_0[3]),.OUT_OBUF(m1_m0_outsel[3]));

	OBUF QL_INST_F2A_B_6_9 (.IN_OBUF(m1_m0_outsel_dup_0[2]),.OUT_OBUF(m1_m0_outsel[2]));

	OBUF QL_INST_F2A_B_6_10 (.IN_OBUF(m1_m0_outsel_dup_0[1]),.OUT_OBUF(m1_m0_outsel[1]));

	OBUF QL_INST_F2A_B_6_11 (.IN_OBUF(m1_m0_outsel_dup_0[0]),.OUT_OBUF(m1_m0_outsel[0]));

	OBUF QL_INST_F2A_B_6_12 (.IN_OBUF(m1_m0_sat_dup_0),.OUT_OBUF(m1_m0_sat));

	OBUF QL_INST_F2A_B_6_13 (.IN_OBUF(m1_m0_rnd_dup_0),.OUT_OBUF(m1_m0_rnd));

	OBUF QL_INST_F2A_B_6_14 (.IN_OBUF(m1_m0_clr_dup_0),.OUT_OBUF(m1_m0_clr));

	OBUF QL_INST_F2A_B_6_15 (.IN_OBUF(m1_oper0_rdata_int[31]),.OUT_OBUF(m1_m0_oper_in[31]));

	OBUF QL_INST_F2A_B_6_16 (.IN_OBUF(m1_oper0_rdata_int[30]),.OUT_OBUF(m1_m0_oper_in[30]));

	OBUF QL_INST_F2A_B_6_17 (.IN_OBUF(m1_oper0_rdata_int[29]),.OUT_OBUF(m1_m0_oper_in[29]));

	DBUF QL_INST_F2Adef_B_6_1 (.IN_DBUF(GND),.OUT_DBUF(m1_oper0_powerdn));

	IBUF QL_INST_A2F_B_6_0 (.IN_IBUF(m1_oper0_rdata[7]),.OUT_IBUF(m1_oper0_rdata_int[7]));

	IBUF QL_INST_A2F_B_6_1 (.IN_IBUF(m1_oper0_rdata[6]),.OUT_IBUF(m1_oper0_rdata_int[6]));

	IBUF QL_INST_A2F_B_6_2 (.IN_IBUF(m1_oper0_rdata[5]),.OUT_IBUF(m1_oper0_rdata_int[5]));

	IBUF QL_INST_A2F_B_6_3 (.IN_IBUF(m1_oper0_rdata[4]),.OUT_IBUF(m1_oper0_rdata_int[4]));

	IBUF QL_INST_A2F_B_6_4 (.IN_IBUF(m1_oper0_rdata[3]),.OUT_IBUF(m1_oper0_rdata_int[3]));

	IBUF QL_INST_A2F_B_6_5 (.IN_IBUF(m1_oper0_rdata[2]),.OUT_IBUF(m1_oper0_rdata_int[2]));

	IBUF QL_INST_A2F_B_6_6 (.IN_IBUF(m1_oper0_rdata[1]),.OUT_IBUF(m1_oper0_rdata_int[1]));

	IBUF QL_INST_A2F_B_6_7 (.IN_IBUF(m1_oper0_rdata[0]),.OUT_IBUF(m1_oper0_rdata_int[0]));

	OBUF QL_INST_F2A_B_7_0 (.IN_OBUF(CLK_int_0__CAND0_BLSBL_7_padClk),.OUT_OBUF(m1_m0_clk));

	OBUF QL_INST_F2A_B_7_1 (.IN_OBUF(m1_oper0_rdata_int[28]),.OUT_OBUF(m1_m0_oper_in[28]));

	OBUF QL_INST_F2A_B_7_2 (.IN_OBUF(m1_oper0_rdata_int[27]),.OUT_OBUF(m1_m0_oper_in[27]));

	OBUF QL_INST_F2A_B_7_3 (.IN_OBUF(m1_oper0_rdata_int[26]),.OUT_OBUF(m1_m0_oper_in[26]));

	OBUF QL_INST_F2A_B_7_4 (.IN_OBUF(m1_oper0_rdata_int[25]),.OUT_OBUF(m1_m0_oper_in[25]));

	OBUF QL_INST_F2A_B_7_5 (.IN_OBUF(m1_oper0_rdata_int[24]),.OUT_OBUF(m1_m0_oper_in[24]));

	OBUF QL_INST_F2A_B_7_6 (.IN_OBUF(m1_oper0_rdata_int[23]),.OUT_OBUF(m1_m0_oper_in[23]));

	OBUF QL_INST_F2A_B_7_7 (.IN_OBUF(m1_oper0_rdata_int[22]),.OUT_OBUF(m1_m0_oper_in[22]));

	OBUF QL_INST_F2A_B_7_8 (.IN_OBUF(m1_oper0_rdata_int[21]),.OUT_OBUF(m1_m0_oper_in[21]));

	OBUF QL_INST_F2A_B_7_9 (.IN_OBUF(m1_oper0_rdata_int[20]),.OUT_OBUF(m1_m0_oper_in[20]));

	OBUF QL_INST_F2A_B_7_10 (.IN_OBUF(m1_oper0_rdata_int[19]),.OUT_OBUF(m1_m0_oper_in[19]));

	OBUF QL_INST_F2A_B_7_11 (.IN_OBUF(m1_oper0_rdata_int[18]),.OUT_OBUF(m1_m0_oper_in[18]));

	IBUF QL_INST_A2F_B_7_0 (.IN_IBUF(m1_m0_dataout[31]),.OUT_IBUF(m1_m0_dataout_int[31]));

	IBUF QL_INST_A2F_B_7_1 (.IN_IBUF(m1_m0_dataout[30]),.OUT_IBUF(m1_m0_dataout_int[30]));

	IBUF QL_INST_A2F_B_7_2 (.IN_IBUF(m1_m0_dataout[29]),.OUT_IBUF(m1_m0_dataout_int[29]));

	IBUF QL_INST_A2F_B_7_3 (.IN_IBUF(m1_m0_dataout[28]),.OUT_IBUF(m1_m0_dataout_int[28]));

	IBUF QL_INST_A2F_B_7_4 (.IN_IBUF(m1_m0_dataout[27]),.OUT_IBUF(m1_m0_dataout_int[27]));

	IBUF QL_INST_A2F_B_7_5 (.IN_IBUF(m1_m0_dataout[26]),.OUT_IBUF(m1_m0_dataout_int[26]));

	OBUF QL_INST_F2A_B_8_0 (.IN_OBUF(m1_oper0_rdata_int[17]),.OUT_OBUF(m1_m0_oper_in[17]));

	OBUF QL_INST_F2A_B_8_1 (.IN_OBUF(m1_oper0_rdata_int[16]),.OUT_OBUF(m1_m0_oper_in[16]));

	OBUF QL_INST_F2A_B_8_2 (.IN_OBUF(m1_oper0_rdata_int[15]),.OUT_OBUF(m1_m0_oper_in[15]));

	OBUF QL_INST_F2A_B_8_3 (.IN_OBUF(m1_oper0_rdata_int[14]),.OUT_OBUF(m1_m0_oper_in[14]));

	OBUF QL_INST_F2A_B_8_4 (.IN_OBUF(m1_oper0_rdata_int[13]),.OUT_OBUF(m1_m0_oper_in[13]));

	OBUF QL_INST_F2A_B_8_5 (.IN_OBUF(m1_oper0_rdata_int[12]),.OUT_OBUF(m1_m0_oper_in[12]));

	OBUF QL_INST_F2A_B_8_6 (.IN_OBUF(m1_oper0_rdata_int[11]),.OUT_OBUF(m1_m0_oper_in[11]));

	OBUF QL_INST_F2A_B_8_7 (.IN_OBUF(m1_oper0_rdata_int[10]),.OUT_OBUF(m1_m0_oper_in[10]));

	OBUF QL_INST_F2A_B_8_8 (.IN_OBUF(m1_oper0_rdata_int[9]),.OUT_OBUF(m1_m0_oper_in[9]));

	OBUF QL_INST_F2A_B_8_9 (.IN_OBUF(m1_oper0_rdata_int[8]),.OUT_OBUF(m1_m0_oper_in[8]));

	OBUF QL_INST_F2A_B_8_10 (.IN_OBUF(m1_oper0_rdata_int[7]),.OUT_OBUF(m1_m0_oper_in[7]));

	OBUF QL_INST_F2A_B_8_11 (.IN_OBUF(m1_oper0_rdata_int[6]),.OUT_OBUF(m1_m0_oper_in[6]));

	OBUF QL_INST_F2A_B_8_12 (.IN_OBUF(m1_oper0_rdata_int[5]),.OUT_OBUF(m1_m0_oper_in[5]));

	OBUF QL_INST_F2A_B_8_13 (.IN_OBUF(m1_oper0_rdata_int[4]),.OUT_OBUF(m1_m0_oper_in[4]));

	OBUF QL_INST_F2A_B_8_14 (.IN_OBUF(m1_oper0_rdata_int[3]),.OUT_OBUF(m1_m0_oper_in[3]));

	OBUF QL_INST_F2A_B_8_15 (.IN_OBUF(m1_oper0_rdata_int[2]),.OUT_OBUF(m1_m0_oper_in[2]));

	OBUF QL_INST_F2A_B_8_16 (.IN_OBUF(m1_oper0_rdata_int[1]),.OUT_OBUF(m1_m0_oper_in[1]));

	OBUF QL_INST_F2A_B_8_17 (.IN_OBUF(m1_oper0_rdata_int[0]),.OUT_OBUF(m1_m0_oper_in[0]));

	IBUF QL_INST_A2F_B_8_0 (.IN_IBUF(m1_m0_dataout[25]),.OUT_IBUF(m1_m0_dataout_int[25]));

	IBUF QL_INST_A2F_B_8_1 (.IN_IBUF(m1_m0_dataout[24]),.OUT_IBUF(m1_m0_dataout_int[24]));

	IBUF QL_INST_A2F_B_8_2 (.IN_IBUF(m1_m0_dataout[23]),.OUT_IBUF(m1_m0_dataout_int[23]));

	IBUF QL_INST_A2F_B_8_3 (.IN_IBUF(m1_m0_dataout[22]),.OUT_IBUF(m1_m0_dataout_int[22]));

	IBUF QL_INST_A2F_B_8_4 (.IN_IBUF(m1_m0_dataout[21]),.OUT_IBUF(m1_m0_dataout_int[21]));

	IBUF QL_INST_A2F_B_8_5 (.IN_IBUF(m1_m0_dataout[20]),.OUT_IBUF(m1_m0_dataout_int[20]));

	IBUF QL_INST_A2F_B_8_6 (.IN_IBUF(m1_m0_dataout[19]),.OUT_IBUF(m1_m0_dataout_int[19]));

	IBUF QL_INST_A2F_B_8_7 (.IN_IBUF(m1_m0_dataout[18]),.OUT_IBUF(m1_m0_dataout_int[18]));

	OBUF QL_INST_F2A_B_9_0 (.IN_OBUF(m1_m0_csel_dup_0),.OUT_OBUF(m1_m0_csel));

	OBUF QL_INST_F2A_B_9_1 (.IN_OBUF(m1_coef_rdata_int[31]),.OUT_OBUF(m1_m0_coef_in[31]));

	OBUF QL_INST_F2A_B_9_2 (.IN_OBUF(m1_coef_rdata_int[30]),.OUT_OBUF(m1_m0_coef_in[30]));

	OBUF QL_INST_F2A_B_9_3 (.IN_OBUF(m1_coef_rdata_int[29]),.OUT_OBUF(m1_m0_coef_in[29]));

	OBUF QL_INST_F2A_B_9_4 (.IN_OBUF(m1_coef_rdata_int[28]),.OUT_OBUF(m1_m0_coef_in[28]));

	OBUF QL_INST_F2A_B_9_5 (.IN_OBUF(m1_coef_rdata_int[27]),.OUT_OBUF(m1_m0_coef_in[27]));

	OBUF QL_INST_F2A_B_9_6 (.IN_OBUF(m1_coef_rdata_int[26]),.OUT_OBUF(m1_m0_coef_in[26]));

	OBUF QL_INST_F2A_B_9_7 (.IN_OBUF(m1_coef_rdata_int[25]),.OUT_OBUF(m1_m0_coef_in[25]));

	OBUF QL_INST_F2A_B_9_8 (.IN_OBUF(m1_coef_rdata_int[24]),.OUT_OBUF(m1_m0_coef_in[24]));

	OBUF QL_INST_F2A_B_9_9 (.IN_OBUF(m1_coef_rdata_int[23]),.OUT_OBUF(m1_m0_coef_in[23]));

	OBUF QL_INST_F2A_B_9_10 (.IN_OBUF(m1_coef_rdata_int[22]),.OUT_OBUF(m1_m0_coef_in[22]));

	OBUF QL_INST_F2A_B_9_11 (.IN_OBUF(m1_coef_rdata_int[21]),.OUT_OBUF(m1_m0_coef_in[21]));

	IBUF QL_INST_A2F_B_9_0 (.IN_IBUF(m1_m0_dataout[17]),.OUT_IBUF(m1_m0_dataout_int[17]));

	IBUF QL_INST_A2F_B_9_1 (.IN_IBUF(m1_m0_dataout[16]),.OUT_IBUF(m1_m0_dataout_int[16]));

	IBUF QL_INST_A2F_B_9_2 (.IN_IBUF(m1_m0_dataout[15]),.OUT_IBUF(m1_m0_dataout_int[15]));

	IBUF QL_INST_A2F_B_9_3 (.IN_IBUF(m1_m0_dataout[14]),.OUT_IBUF(m1_m0_dataout_int[14]));

	IBUF QL_INST_A2F_B_9_4 (.IN_IBUF(m1_m0_dataout[13]),.OUT_IBUF(m1_m0_dataout_int[13]));

	IBUF QL_INST_A2F_B_9_5 (.IN_IBUF(m1_m0_dataout[12]),.OUT_IBUF(m1_m0_dataout_int[12]));

	OBUF QL_INST_F2A_B_10_0 (.IN_OBUF(m1_coef_rdata_int[20]),.OUT_OBUF(m1_m0_coef_in[20]));

	OBUF QL_INST_F2A_B_10_1 (.IN_OBUF(m1_coef_rdata_int[19]),.OUT_OBUF(m1_m0_coef_in[19]));

	OBUF QL_INST_F2A_B_10_2 (.IN_OBUF(m1_coef_rdata_int[18]),.OUT_OBUF(m1_m0_coef_in[18]));

	OBUF QL_INST_F2A_B_10_3 (.IN_OBUF(m1_coef_rdata_int[17]),.OUT_OBUF(m1_m0_coef_in[17]));

	OBUF QL_INST_F2A_B_10_4 (.IN_OBUF(m1_coef_rdata_int[16]),.OUT_OBUF(m1_m0_coef_in[16]));

	OBUF QL_INST_F2A_B_10_5 (.IN_OBUF(m1_coef_rdata_int[15]),.OUT_OBUF(m1_m0_coef_in[15]));

	OBUF QL_INST_F2A_B_10_6 (.IN_OBUF(m1_coef_rdata_int[14]),.OUT_OBUF(m1_m0_coef_in[14]));

	OBUF QL_INST_F2A_B_10_7 (.IN_OBUF(m1_coef_rdata_int[13]),.OUT_OBUF(m1_m0_coef_in[13]));

	OBUF QL_INST_F2A_B_10_8 (.IN_OBUF(m1_coef_rdata_int[12]),.OUT_OBUF(m1_m0_coef_in[12]));

	OBUF QL_INST_F2A_B_10_9 (.IN_OBUF(m1_coef_rdata_int[11]),.OUT_OBUF(m1_m0_coef_in[11]));

	OBUF QL_INST_F2A_B_10_10 (.IN_OBUF(m1_coef_rdata_int[10]),.OUT_OBUF(m1_m0_coef_in[10]));

	OBUF QL_INST_F2A_B_10_11 (.IN_OBUF(m1_coef_rdata_int[9]),.OUT_OBUF(m1_m0_coef_in[9]));

	OBUF QL_INST_F2A_B_10_12 (.IN_OBUF(m1_coef_rdata_int[8]),.OUT_OBUF(m1_m0_coef_in[8]));

	OBUF QL_INST_F2A_B_10_13 (.IN_OBUF(m1_coef_rdata_int[7]),.OUT_OBUF(m1_m0_coef_in[7]));

	OBUF QL_INST_F2A_B_10_14 (.IN_OBUF(m1_coef_rdata_int[6]),.OUT_OBUF(m1_m0_coef_in[6]));

	OBUF QL_INST_F2A_B_10_15 (.IN_OBUF(m1_coef_rdata_int[5]),.OUT_OBUF(m1_m0_coef_in[5]));

	OBUF QL_INST_F2A_B_10_16 (.IN_OBUF(m1_coef_rdata_int[4]),.OUT_OBUF(m1_m0_coef_in[4]));

	OBUF QL_INST_F2A_B_10_17 (.IN_OBUF(m1_coef_rdata_int[3]),.OUT_OBUF(m1_m0_coef_in[3]));

	IBUF QL_INST_A2F_B_10_0 (.IN_IBUF(m1_m0_dataout[11]),.OUT_IBUF(m1_m0_dataout_int[11]));

	IBUF QL_INST_A2F_B_10_1 (.IN_IBUF(m1_m0_dataout[10]),.OUT_IBUF(m1_m0_dataout_int[10]));

	IBUF QL_INST_A2F_B_10_2 (.IN_IBUF(m1_m0_dataout[9]),.OUT_IBUF(m1_m0_dataout_int[9]));

	IBUF QL_INST_A2F_B_10_3 (.IN_IBUF(m1_m0_dataout[8]),.OUT_IBUF(m1_m0_dataout_int[8]));

	IBUF QL_INST_A2F_B_10_4 (.IN_IBUF(m1_m0_dataout[7]),.OUT_IBUF(m1_m0_dataout_int[7]));

	IBUF QL_INST_A2F_B_10_5 (.IN_IBUF(m1_m0_dataout[6]),.OUT_IBUF(m1_m0_dataout_int[6]));

	IBUF QL_INST_A2F_B_10_6 (.IN_IBUF(m1_m0_dataout[5]),.OUT_IBUF(m1_m0_dataout_int[5]));

	IBUF QL_INST_A2F_B_10_7 (.IN_IBUF(m1_m0_dataout[4]),.OUT_IBUF(m1_m0_dataout_int[4]));

	OBUF QL_INST_F2A_B_11_0 (.IN_OBUF(m1_coef_rdata_int[2]),.OUT_OBUF(m1_m0_coef_in[2]));

	OBUF QL_INST_F2A_B_11_1 (.IN_OBUF(m1_coef_rdata_int[1]),.OUT_OBUF(m1_m0_coef_in[1]));

	OBUF QL_INST_F2A_B_11_2 (.IN_OBUF(m1_coef_rdata_int[0]),.OUT_OBUF(m1_m0_coef_in[0]));

	OBUF QL_INST_F2A_B_11_3 (.IN_OBUF(m1_m0_mode_dup_0[1]),.OUT_OBUF(m1_m0_mode[1]));

	OBUF QL_INST_F2A_B_11_4 (.IN_OBUF(m1_m0_mode_dup_0[0]),.OUT_OBUF(m1_m0_mode[0]));

	OBUF QL_INST_F2A_B_11_5 (.IN_OBUF(m1_m0_tc_dup_0),.OUT_OBUF(m1_m0_tc));

	OBUF QL_INST_F2A_B_11_6 (.IN_OBUF(m1_m0_reset_dup_0),.OUT_OBUF(m1_m0_reset));

	OBUF QL_INST_F2A_B_11_7 (.IN_OBUF(m1_coef_wdata_dup_0[31]),.OUT_OBUF(m1_coef_wdata[31]));

	OBUF QL_INST_F2A_B_11_8 (.IN_OBUF(m1_coef_wdata_dup_0[30]),.OUT_OBUF(m1_coef_wdata[30]));

	OBUF QL_INST_F2A_B_11_9 (.IN_OBUF(m1_coef_wdata_dup_0[29]),.OUT_OBUF(m1_coef_wdata[29]));

	OBUF QL_INST_F2A_B_11_10 (.IN_OBUF(m1_coef_wdata_dup_0[28]),.OUT_OBUF(m1_coef_wdata[28]));

	OBUF QL_INST_F2A_B_11_11 (.IN_OBUF(m1_coef_wdata_dup_0[27]),.OUT_OBUF(m1_coef_wdata[27]));

	IBUF QL_INST_A2F_B_11_0 (.IN_IBUF(m1_m0_dataout[3]),.OUT_IBUF(m1_m0_dataout_int[3]));

	IBUF QL_INST_A2F_B_11_1 (.IN_IBUF(m1_m0_dataout[2]),.OUT_IBUF(m1_m0_dataout_int[2]));

	IBUF QL_INST_A2F_B_11_2 (.IN_IBUF(m1_m0_dataout[1]),.OUT_IBUF(m1_m0_dataout_int[1]));

	IBUF QL_INST_A2F_B_11_3 (.IN_IBUF(m1_m0_dataout[0]),.OUT_IBUF(m1_m0_dataout_int[0]));

	IBUF QL_INST_A2F_B_11_4 (.IN_IBUF(m1_coef_rdata[31]),.OUT_IBUF(m1_coef_rdata_int[31]));

	IBUF QL_INST_A2F_B_11_5 (.IN_IBUF(m1_coef_rdata[30]),.OUT_IBUF(m1_coef_rdata_int[30]));

	OBUF QL_INST_F2A_B_12_0 (.IN_OBUF(m1_coef_wdata_dup_0[26]),.OUT_OBUF(m1_coef_wdata[26]));

	OBUF QL_INST_F2A_B_12_1 (.IN_OBUF(m1_coef_wdata_dup_0[25]),.OUT_OBUF(m1_coef_wdata[25]));

	OBUF QL_INST_F2A_B_12_2 (.IN_OBUF(m1_coef_wdata_dup_0[24]),.OUT_OBUF(m1_coef_wdata[24]));

	OBUF QL_INST_F2A_B_12_3 (.IN_OBUF(m1_coef_wdata_dup_0[23]),.OUT_OBUF(m1_coef_wdata[23]));

	OBUF QL_INST_F2A_B_12_4 (.IN_OBUF(m1_coef_wdata_dup_0[22]),.OUT_OBUF(m1_coef_wdata[22]));

	OBUF QL_INST_F2A_B_12_5 (.IN_OBUF(m1_coef_wdata_dup_0[21]),.OUT_OBUF(m1_coef_wdata[21]));

	OBUF QL_INST_F2A_B_12_6 (.IN_OBUF(m1_coef_wdata_dup_0[20]),.OUT_OBUF(m1_coef_wdata[20]));

	OBUF QL_INST_F2A_B_12_7 (.IN_OBUF(m1_coef_wdata_dup_0[19]),.OUT_OBUF(m1_coef_wdata[19]));

	OBUF QL_INST_F2A_B_12_8 (.IN_OBUF(m1_coef_wdata_dup_0[18]),.OUT_OBUF(m1_coef_wdata[18]));

	OBUF QL_INST_F2A_B_12_9 (.IN_OBUF(m1_coef_wdata_dup_0[17]),.OUT_OBUF(m1_coef_wdata[17]));

	OBUF QL_INST_F2A_B_12_10 (.IN_OBUF(m1_coef_wdata_dup_0[16]),.OUT_OBUF(m1_coef_wdata[16]));

	OBUF QL_INST_F2A_B_12_11 (.IN_OBUF(m1_coef_wdata_dup_0[15]),.OUT_OBUF(m1_coef_wdata[15]));

	OBUF QL_INST_F2A_B_12_12 (.IN_OBUF(m1_coef_wdata_dup_0[14]),.OUT_OBUF(m1_coef_wdata[14]));

	OBUF QL_INST_F2A_B_12_13 (.IN_OBUF(m1_coef_wdata_dup_0[13]),.OUT_OBUF(m1_coef_wdata[13]));

	OBUF QL_INST_F2A_B_12_14 (.IN_OBUF(m1_coef_wdata_dup_0[12]),.OUT_OBUF(m1_coef_wdata[12]));

	OBUF QL_INST_F2A_B_12_15 (.IN_OBUF(m1_coef_wdata_dup_0[11]),.OUT_OBUF(m1_coef_wdata[11]));

	OBUF QL_INST_F2A_B_12_16 (.IN_OBUF(m1_coef_wdata_dup_0[10]),.OUT_OBUF(m1_coef_wdata[10]));

	OBUF QL_INST_F2A_B_12_17 (.IN_OBUF(m1_coef_wdata_dup_0[9]),.OUT_OBUF(m1_coef_wdata[9]));

	IBUF QL_INST_A2F_B_12_0 (.IN_IBUF(m1_coef_rdata[29]),.OUT_IBUF(m1_coef_rdata_int[29]));

	IBUF QL_INST_A2F_B_12_1 (.IN_IBUF(m1_coef_rdata[28]),.OUT_IBUF(m1_coef_rdata_int[28]));

	IBUF QL_INST_A2F_B_12_2 (.IN_IBUF(m1_coef_rdata[27]),.OUT_IBUF(m1_coef_rdata_int[27]));

	IBUF QL_INST_A2F_B_12_3 (.IN_IBUF(m1_coef_rdata[26]),.OUT_IBUF(m1_coef_rdata_int[26]));

	IBUF QL_INST_A2F_B_12_4 (.IN_IBUF(m1_coef_rdata[25]),.OUT_IBUF(m1_coef_rdata_int[25]));

	IBUF QL_INST_A2F_B_12_5 (.IN_IBUF(m1_coef_rdata[24]),.OUT_IBUF(m1_coef_rdata_int[24]));

	IBUF QL_INST_A2F_B_12_6 (.IN_IBUF(m1_coef_rdata[23]),.OUT_IBUF(m1_coef_rdata_int[23]));

	IBUF QL_INST_A2F_B_12_7 (.IN_IBUF(m1_coef_rdata[22]),.OUT_IBUF(m1_coef_rdata_int[22]));

	OBUF QL_INST_F2A_B_13_0 (.IN_OBUF(CLK_int_0__CAND0_BLSBR_13_padClk),.OUT_OBUF(m1_coef_wclk));

	OBUF QL_INST_F2A_B_13_1 (.IN_OBUF(m1_coef_wdata_dup_0[8]),.OUT_OBUF(m1_coef_wdata[8]));

	OBUF QL_INST_F2A_B_13_2 (.IN_OBUF(m1_coef_wdata_dup_0[7]),.OUT_OBUF(m1_coef_wdata[7]));

	OBUF QL_INST_F2A_B_13_3 (.IN_OBUF(m1_coef_wdata_dup_0[6]),.OUT_OBUF(m1_coef_wdata[6]));

	OBUF QL_INST_F2A_B_13_4 (.IN_OBUF(m1_coef_wdata_dup_0[5]),.OUT_OBUF(m1_coef_wdata[5]));

	OBUF QL_INST_F2A_B_13_5 (.IN_OBUF(m1_coef_wdata_dup_0[4]),.OUT_OBUF(m1_coef_wdata[4]));

	OBUF QL_INST_F2A_B_13_6 (.IN_OBUF(m1_coef_wdata_dup_0[3]),.OUT_OBUF(m1_coef_wdata[3]));

	OBUF QL_INST_F2A_B_13_7 (.IN_OBUF(m1_coef_wdata_dup_0[2]),.OUT_OBUF(m1_coef_wdata[2]));

	OBUF QL_INST_F2A_B_13_8 (.IN_OBUF(m1_coef_wdata_dup_0[1]),.OUT_OBUF(m1_coef_wdata[1]));

	OBUF QL_INST_F2A_B_13_9 (.IN_OBUF(m1_coef_wdata_dup_0[0]),.OUT_OBUF(m1_coef_wdata[0]));

	OBUF QL_INST_F2A_B_13_10 (.IN_OBUF(m1_coef_waddr_dup_0[11]),.OUT_OBUF(m1_coef_waddr[11]));

	OBUF QL_INST_F2A_B_13_11 (.IN_OBUF(m1_coef_waddr_dup_0[10]),.OUT_OBUF(m1_coef_waddr[10]));

	DBUF QL_INST_F2Adef_B_13_0 (.IN_DBUF(GND),.OUT_DBUF(m1_coef_powerdn));

	IBUF QL_INST_A2F_B_13_0 (.IN_IBUF(m1_coef_rdata[21]),.OUT_IBUF(m1_coef_rdata_int[21]));

	IBUF QL_INST_A2F_B_13_1 (.IN_IBUF(m1_coef_rdata[20]),.OUT_IBUF(m1_coef_rdata_int[20]));

	IBUF QL_INST_A2F_B_13_2 (.IN_IBUF(m1_coef_rdata[19]),.OUT_IBUF(m1_coef_rdata_int[19]));

	IBUF QL_INST_A2F_B_13_3 (.IN_IBUF(m1_coef_rdata[18]),.OUT_IBUF(m1_coef_rdata_int[18]));

	IBUF QL_INST_A2F_B_13_4 (.IN_IBUF(m1_coef_rdata[17]),.OUT_IBUF(m1_coef_rdata_int[17]));

	IBUF QL_INST_A2F_B_13_5 (.IN_IBUF(m1_coef_rdata[16]),.OUT_IBUF(m1_coef_rdata_int[16]));

	OBUF QL_INST_F2A_B_14_0 (.IN_OBUF(m1_coef_waddr_dup_0[9]),.OUT_OBUF(m1_coef_waddr[9]));

	OBUF QL_INST_F2A_B_14_1 (.IN_OBUF(m1_coef_waddr_dup_0[8]),.OUT_OBUF(m1_coef_waddr[8]));

	OBUF QL_INST_F2A_B_14_2 (.IN_OBUF(m1_coef_waddr_dup_0[7]),.OUT_OBUF(m1_coef_waddr[7]));

	OBUF QL_INST_F2A_B_14_3 (.IN_OBUF(m1_coef_waddr_dup_0[6]),.OUT_OBUF(m1_coef_waddr[6]));

	OBUF QL_INST_F2A_B_14_4 (.IN_OBUF(m1_coef_waddr_dup_0[5]),.OUT_OBUF(m1_coef_waddr[5]));

	OBUF QL_INST_F2A_B_14_5 (.IN_OBUF(m1_coef_waddr_dup_0[4]),.OUT_OBUF(m1_coef_waddr[4]));

	OBUF QL_INST_F2A_B_14_6 (.IN_OBUF(m1_coef_waddr_dup_0[3]),.OUT_OBUF(m1_coef_waddr[3]));

	OBUF QL_INST_F2A_B_14_7 (.IN_OBUF(m1_coef_waddr_dup_0[2]),.OUT_OBUF(m1_coef_waddr[2]));

	OBUF QL_INST_F2A_B_14_8 (.IN_OBUF(m1_coef_waddr_dup_0[1]),.OUT_OBUF(m1_coef_waddr[1]));

	OBUF QL_INST_F2A_B_14_9 (.IN_OBUF(m1_coef_waddr_dup_0[0]),.OUT_OBUF(m1_coef_waddr[0]));

	OBUF QL_INST_F2A_B_14_10 (.IN_OBUF(m1_coef_we_dup_0),.OUT_OBUF(m1_coef_we));

	OBUF QL_INST_F2A_B_14_11 (.IN_OBUF(m0_coef_wdsel_dup_0),.OUT_OBUF(m1_coef_wdsel));

	OBUF QL_INST_F2A_B_14_12 (.IN_OBUF(m0_coef_rmode_dup_0[1]),.OUT_OBUF(m1_coef_rmode[1]));

	OBUF QL_INST_F2A_B_14_13 (.IN_OBUF(m0_coef_rmode_dup_0[0]),.OUT_OBUF(m1_coef_rmode[0]));

	OBUF QL_INST_F2A_B_14_14 (.IN_OBUF(m1_coef_raddr_dup_0[11]),.OUT_OBUF(m1_coef_raddr[11]));

	OBUF QL_INST_F2A_B_14_15 (.IN_OBUF(m1_coef_raddr_dup_0[10]),.OUT_OBUF(m1_coef_raddr[10]));

	OBUF QL_INST_F2A_B_14_16 (.IN_OBUF(m1_coef_raddr_dup_0[9]),.OUT_OBUF(m1_coef_raddr[9]));

	OBUF QL_INST_F2A_B_14_17 (.IN_OBUF(m1_coef_raddr_dup_0[8]),.OUT_OBUF(m1_coef_raddr[8]));

	IBUF QL_INST_A2F_B_14_0 (.IN_IBUF(m1_coef_rdata[15]),.OUT_IBUF(m1_coef_rdata_int[15]));

	IBUF QL_INST_A2F_B_14_1 (.IN_IBUF(m1_coef_rdata[14]),.OUT_IBUF(m1_coef_rdata_int[14]));

	IBUF QL_INST_A2F_B_14_2 (.IN_IBUF(m1_coef_rdata[13]),.OUT_IBUF(m1_coef_rdata_int[13]));

	IBUF QL_INST_A2F_B_14_3 (.IN_IBUF(m1_coef_rdata[12]),.OUT_IBUF(m1_coef_rdata_int[12]));

	IBUF QL_INST_A2F_B_14_4 (.IN_IBUF(m1_coef_rdata[11]),.OUT_IBUF(m1_coef_rdata_int[11]));

	IBUF QL_INST_A2F_B_14_5 (.IN_IBUF(m1_coef_rdata[10]),.OUT_IBUF(m1_coef_rdata_int[10]));

	IBUF QL_INST_A2F_B_14_6 (.IN_IBUF(m1_coef_rdata[9]),.OUT_IBUF(m1_coef_rdata_int[9]));

	IBUF QL_INST_A2F_B_14_7 (.IN_IBUF(m1_coef_rdata[8]),.OUT_IBUF(m1_coef_rdata_int[8]));

	OBUF QL_INST_F2A_B_15_0 (.IN_OBUF(CLK_int_0__CAND0_BLSBR_15_padClk),.OUT_OBUF(m1_coef_rclk));

	OBUF QL_INST_F2A_B_15_1 (.IN_OBUF(m1_coef_raddr_dup_0[7]),.OUT_OBUF(m1_coef_raddr[7]));

	OBUF QL_INST_F2A_B_15_2 (.IN_OBUF(m1_coef_raddr_dup_0[6]),.OUT_OBUF(m1_coef_raddr[6]));

	OBUF QL_INST_F2A_B_15_3 (.IN_OBUF(m1_coef_raddr_dup_0[5]),.OUT_OBUF(m1_coef_raddr[5]));

	OBUF QL_INST_F2A_B_15_4 (.IN_OBUF(m1_coef_raddr_dup_0[4]),.OUT_OBUF(m1_coef_raddr[4]));

	OBUF QL_INST_F2A_B_15_5 (.IN_OBUF(m1_coef_raddr_dup_0[3]),.OUT_OBUF(m1_coef_raddr[3]));

	OBUF QL_INST_F2A_B_15_6 (.IN_OBUF(m1_coef_raddr_dup_0[2]),.OUT_OBUF(m1_coef_raddr[2]));

	OBUF QL_INST_F2A_B_15_7 (.IN_OBUF(m1_coef_raddr_dup_0[1]),.OUT_OBUF(m1_coef_raddr[1]));

	OBUF QL_INST_F2A_B_15_8 (.IN_OBUF(m1_coef_raddr_dup_0[0]),.OUT_OBUF(m1_coef_raddr[0]));

	OBUF QL_INST_F2A_B_15_9 (.IN_OBUF(m0_coef_wmode_dup_0[1]),.OUT_OBUF(m1_coef_wmode[1]));

	OBUF QL_INST_F2A_B_15_10 (.IN_OBUF(m0_coef_wmode_dup_0[0]),.OUT_OBUF(m1_coef_wmode[0]));

	IBUF QL_INST_A2F_B_15_0 (.IN_IBUF(m1_coef_rdata[7]),.OUT_IBUF(m1_coef_rdata_int[7]));

	IBUF QL_INST_A2F_B_15_1 (.IN_IBUF(m1_coef_rdata[6]),.OUT_IBUF(m1_coef_rdata_int[6]));

	IBUF QL_INST_A2F_B_15_2 (.IN_IBUF(m1_coef_rdata[5]),.OUT_IBUF(m1_coef_rdata_int[5]));

	IBUF QL_INST_A2F_B_15_3 (.IN_IBUF(m1_coef_rdata[4]),.OUT_IBUF(m1_coef_rdata_int[4]));

	IBUF QL_INST_A2F_B_15_4 (.IN_IBUF(m1_coef_rdata[3]),.OUT_IBUF(m1_coef_rdata_int[3]));

	IBUF QL_INST_A2F_B_15_5 (.IN_IBUF(m1_coef_rdata[2]),.OUT_IBUF(m1_coef_rdata_int[2]));

	IBUF QL_INST_A2F_B_16_0 (.IN_IBUF(m1_coef_rdata[1]),.OUT_IBUF(m1_coef_rdata_int[1]));

	IBUF QL_INST_A2F_B_16_1 (.IN_IBUF(m1_coef_rdata[0]),.OUT_IBUF(m1_coef_rdata_int[0]));

	OBUF QL_INST_F2A_B_18_7 (.IN_OBUF(m0_m0_outsel_dup_0[5]),.OUT_OBUF(m1_m1_outsel[5]));

	OBUF QL_INST_F2A_B_18_8 (.IN_OBUF(m0_m0_outsel_dup_0[4]),.OUT_OBUF(m1_m1_outsel[4]));

	OBUF QL_INST_F2A_B_18_9 (.IN_OBUF(m0_m0_outsel_dup_0[3]),.OUT_OBUF(m1_m1_outsel[3]));

	OBUF QL_INST_F2A_B_18_10 (.IN_OBUF(m0_m0_outsel_dup_0[2]),.OUT_OBUF(m1_m1_outsel[2]));

	OBUF QL_INST_F2A_B_18_11 (.IN_OBUF(m0_m0_outsel_dup_0[1]),.OUT_OBUF(m1_m1_outsel[1]));

	OBUF QL_INST_F2A_B_18_12 (.IN_OBUF(m0_m0_outsel_dup_0[0]),.OUT_OBUF(m1_m1_outsel[0]));

	OBUF QL_INST_F2A_B_18_13 (.IN_OBUF(m1_m1_sat_dup_0),.OUT_OBUF(m1_m1_sat));

	OBUF QL_INST_F2A_B_18_14 (.IN_OBUF(m1_m1_rnd_dup_0),.OUT_OBUF(m1_m1_rnd));

	OBUF QL_INST_F2A_B_18_15 (.IN_OBUF(m1_m1_clr_dup_0),.OUT_OBUF(m1_m1_clr));

	OBUF QL_INST_F2A_B_18_16 (.IN_OBUF(m1_m1_clken_dup_0),.OUT_OBUF(m1_m1_clken));

	IBUF QL_INST_A2F_B_18_6 (.IN_IBUF(m1_m1_dataout[31]),.OUT_IBUF(m1_m1_dataout_int[31]));

	IBUF QL_INST_A2F_B_18_7 (.IN_IBUF(m1_m1_dataout[30]),.OUT_IBUF(m1_m1_dataout_int[30]));

	OBUF QL_INST_F2A_B_19_0 (.IN_OBUF(CLK_int_0__CAND0_BRSBL_19_padClk),.OUT_OBUF(m1_m1_clk));

	OBUF QL_INST_F2A_B_19_1 (.IN_OBUF(m1_m1_osel_dup_0),.OUT_OBUF(m1_m1_osel));

	OBUF QL_INST_F2A_B_19_2 (.IN_OBUF(m1_m1_tc_dup_0),.OUT_OBUF(m1_m1_tc));

	OBUF QL_INST_F2A_B_19_3 (.IN_OBUF(m1_m1_reset_dup_0),.OUT_OBUF(m1_m1_reset));

	OBUF QL_INST_F2A_B_19_4 (.IN_OBUF(m1_coef_rdata_int[31]),.OUT_OBUF(m1_m1_coef_in[31]));

	OBUF QL_INST_F2A_B_19_5 (.IN_OBUF(m1_coef_rdata_int[30]),.OUT_OBUF(m1_m1_coef_in[30]));

	OBUF QL_INST_F2A_B_19_6 (.IN_OBUF(m1_coef_rdata_int[29]),.OUT_OBUF(m1_m1_coef_in[29]));

	OBUF QL_INST_F2A_B_19_7 (.IN_OBUF(m1_coef_rdata_int[28]),.OUT_OBUF(m1_m1_coef_in[28]));

	OBUF QL_INST_F2A_B_19_8 (.IN_OBUF(m1_coef_rdata_int[27]),.OUT_OBUF(m1_m1_coef_in[27]));

	OBUF QL_INST_F2A_B_19_9 (.IN_OBUF(m1_coef_rdata_int[26]),.OUT_OBUF(m1_m1_coef_in[26]));

	OBUF QL_INST_F2A_B_19_10 (.IN_OBUF(m1_coef_rdata_int[25]),.OUT_OBUF(m1_m1_coef_in[25]));

	OBUF QL_INST_F2A_B_19_11 (.IN_OBUF(m1_coef_rdata_int[24]),.OUT_OBUF(m1_m1_coef_in[24]));

	IBUF QL_INST_A2F_B_19_0 (.IN_IBUF(m1_m1_dataout[29]),.OUT_IBUF(m1_m1_dataout_int[29]));

	IBUF QL_INST_A2F_B_19_1 (.IN_IBUF(m1_m1_dataout[28]),.OUT_IBUF(m1_m1_dataout_int[28]));

	IBUF QL_INST_A2F_B_19_2 (.IN_IBUF(m1_m1_dataout[27]),.OUT_IBUF(m1_m1_dataout_int[27]));

	IBUF QL_INST_A2F_B_19_3 (.IN_IBUF(m1_m1_dataout[26]),.OUT_IBUF(m1_m1_dataout_int[26]));

	IBUF QL_INST_A2F_B_19_4 (.IN_IBUF(m1_m1_dataout[25]),.OUT_IBUF(m1_m1_dataout_int[25]));

	IBUF QL_INST_A2F_B_19_5 (.IN_IBUF(m1_m1_dataout[24]),.OUT_IBUF(m1_m1_dataout_int[24]));

	OBUF QL_INST_F2A_B_20_0 (.IN_OBUF(m1_coef_rdata_int[23]),.OUT_OBUF(m1_m1_coef_in[23]));

	OBUF QL_INST_F2A_B_20_1 (.IN_OBUF(m1_coef_rdata_int[22]),.OUT_OBUF(m1_m1_coef_in[22]));

	OBUF QL_INST_F2A_B_20_2 (.IN_OBUF(m1_coef_rdata_int[21]),.OUT_OBUF(m1_m1_coef_in[21]));

	OBUF QL_INST_F2A_B_20_3 (.IN_OBUF(m1_coef_rdata_int[20]),.OUT_OBUF(m1_m1_coef_in[20]));

	OBUF QL_INST_F2A_B_20_4 (.IN_OBUF(m1_coef_rdata_int[19]),.OUT_OBUF(m1_m1_coef_in[19]));

	OBUF QL_INST_F2A_B_20_5 (.IN_OBUF(m1_coef_rdata_int[18]),.OUT_OBUF(m1_m1_coef_in[18]));

	OBUF QL_INST_F2A_B_20_6 (.IN_OBUF(m1_coef_rdata_int[17]),.OUT_OBUF(m1_m1_coef_in[17]));

	OBUF QL_INST_F2A_B_20_7 (.IN_OBUF(m1_coef_rdata_int[16]),.OUT_OBUF(m1_m1_coef_in[16]));

	OBUF QL_INST_F2A_B_20_8 (.IN_OBUF(m1_coef_rdata_int[15]),.OUT_OBUF(m1_m1_coef_in[15]));

	OBUF QL_INST_F2A_B_20_9 (.IN_OBUF(m1_coef_rdata_int[14]),.OUT_OBUF(m1_m1_coef_in[14]));

	OBUF QL_INST_F2A_B_20_10 (.IN_OBUF(m1_coef_rdata_int[13]),.OUT_OBUF(m1_m1_coef_in[13]));

	OBUF QL_INST_F2A_B_20_11 (.IN_OBUF(m1_coef_rdata_int[12]),.OUT_OBUF(m1_m1_coef_in[12]));

	OBUF QL_INST_F2A_B_20_12 (.IN_OBUF(m1_coef_rdata_int[11]),.OUT_OBUF(m1_m1_coef_in[11]));

	OBUF QL_INST_F2A_B_20_13 (.IN_OBUF(m1_coef_rdata_int[10]),.OUT_OBUF(m1_m1_coef_in[10]));

	OBUF QL_INST_F2A_B_20_14 (.IN_OBUF(m1_coef_rdata_int[9]),.OUT_OBUF(m1_m1_coef_in[9]));

	OBUF QL_INST_F2A_B_20_15 (.IN_OBUF(m1_coef_rdata_int[8]),.OUT_OBUF(m1_m1_coef_in[8]));

	OBUF QL_INST_F2A_B_20_16 (.IN_OBUF(m1_coef_rdata_int[7]),.OUT_OBUF(m1_m1_coef_in[7]));

	OBUF QL_INST_F2A_B_20_17 (.IN_OBUF(m1_coef_rdata_int[6]),.OUT_OBUF(m1_m1_coef_in[6]));

	IBUF QL_INST_A2F_B_20_0 (.IN_IBUF(m1_m1_dataout[23]),.OUT_IBUF(m1_m1_dataout_int[23]));

	IBUF QL_INST_A2F_B_20_1 (.IN_IBUF(m1_m1_dataout[22]),.OUT_IBUF(m1_m1_dataout_int[22]));

	IBUF QL_INST_A2F_B_20_2 (.IN_IBUF(m1_m1_dataout[21]),.OUT_IBUF(m1_m1_dataout_int[21]));

	IBUF QL_INST_A2F_B_20_3 (.IN_IBUF(m1_m1_dataout[20]),.OUT_IBUF(m1_m1_dataout_int[20]));

	IBUF QL_INST_A2F_B_20_4 (.IN_IBUF(m1_m1_dataout[19]),.OUT_IBUF(m1_m1_dataout_int[19]));

	IBUF QL_INST_A2F_B_20_5 (.IN_IBUF(m1_m1_dataout[18]),.OUT_IBUF(m1_m1_dataout_int[18]));

	IBUF QL_INST_A2F_B_20_6 (.IN_IBUF(m1_m1_dataout[17]),.OUT_IBUF(m1_m1_dataout_int[17]));

	OBUF QL_INST_F2A_B_21_0 (.IN_OBUF(m1_coef_rdata_int[5]),.OUT_OBUF(m1_m1_coef_in[5]));

	OBUF QL_INST_F2A_B_21_1 (.IN_OBUF(m1_coef_rdata_int[4]),.OUT_OBUF(m1_m1_coef_in[4]));

	OBUF QL_INST_F2A_B_21_2 (.IN_OBUF(m1_coef_rdata_int[3]),.OUT_OBUF(m1_m1_coef_in[3]));

	OBUF QL_INST_F2A_B_21_3 (.IN_OBUF(m1_coef_rdata_int[2]),.OUT_OBUF(m1_m1_coef_in[2]));

	OBUF QL_INST_F2A_B_21_4 (.IN_OBUF(m1_coef_rdata_int[1]),.OUT_OBUF(m1_m1_coef_in[1]));

	OBUF QL_INST_F2A_B_21_5 (.IN_OBUF(m1_coef_rdata_int[0]),.OUT_OBUF(m1_m1_coef_in[0]));

	OBUF QL_INST_F2A_B_21_6 (.IN_OBUF(m1_m1_mode_dup_0[1]),.OUT_OBUF(m1_m1_mode[1]));

	OBUF QL_INST_F2A_B_21_7 (.IN_OBUF(m1_m1_csel_dup_0),.OUT_OBUF(m1_m1_csel));

	OBUF QL_INST_F2A_B_21_8 (.IN_OBUF(m1_m1_mode_dup_0[0]),.OUT_OBUF(m1_m1_mode[0]));

	OBUF QL_INST_F2A_B_21_9 (.IN_OBUF(m1_oper1_rdata_int[31]),.OUT_OBUF(m1_m1_oper_in[31]));

	OBUF QL_INST_F2A_B_21_10 (.IN_OBUF(m1_oper1_rdata_int[30]),.OUT_OBUF(m1_m1_oper_in[30]));

	OBUF QL_INST_F2A_B_21_11 (.IN_OBUF(m1_oper1_rdata_int[29]),.OUT_OBUF(m1_m1_oper_in[29]));

	IBUF QL_INST_A2F_B_21_0 (.IN_IBUF(m1_m1_dataout[16]),.OUT_IBUF(m1_m1_dataout_int[16]));

	IBUF QL_INST_A2F_B_21_1 (.IN_IBUF(m1_m1_dataout[15]),.OUT_IBUF(m1_m1_dataout_int[15]));

	IBUF QL_INST_A2F_B_21_2 (.IN_IBUF(m1_m1_dataout[14]),.OUT_IBUF(m1_m1_dataout_int[14]));

	IBUF QL_INST_A2F_B_21_3 (.IN_IBUF(m1_m1_dataout[13]),.OUT_IBUF(m1_m1_dataout_int[13]));

	IBUF QL_INST_A2F_B_21_4 (.IN_IBUF(m1_m1_dataout[12]),.OUT_IBUF(m1_m1_dataout_int[12]));

	IBUF QL_INST_A2F_B_21_5 (.IN_IBUF(m1_m1_dataout[11]),.OUT_IBUF(m1_m1_dataout_int[11]));

	OBUF QL_INST_F2A_B_22_0 (.IN_OBUF(m1_oper1_rdata_int[28]),.OUT_OBUF(m1_m1_oper_in[28]));

	OBUF QL_INST_F2A_B_22_1 (.IN_OBUF(m1_oper1_rdata_int[27]),.OUT_OBUF(m1_m1_oper_in[27]));

	OBUF QL_INST_F2A_B_22_2 (.IN_OBUF(m1_oper1_rdata_int[26]),.OUT_OBUF(m1_m1_oper_in[26]));

	OBUF QL_INST_F2A_B_22_3 (.IN_OBUF(m1_oper1_rdata_int[25]),.OUT_OBUF(m1_m1_oper_in[25]));

	OBUF QL_INST_F2A_B_22_4 (.IN_OBUF(m1_oper1_rdata_int[24]),.OUT_OBUF(m1_m1_oper_in[24]));

	OBUF QL_INST_F2A_B_22_5 (.IN_OBUF(m1_oper1_rdata_int[23]),.OUT_OBUF(m1_m1_oper_in[23]));

	OBUF QL_INST_F2A_B_22_6 (.IN_OBUF(m1_oper1_rdata_int[22]),.OUT_OBUF(m1_m1_oper_in[22]));

	OBUF QL_INST_F2A_B_22_7 (.IN_OBUF(m1_oper1_rdata_int[21]),.OUT_OBUF(m1_m1_oper_in[21]));

	OBUF QL_INST_F2A_B_22_8 (.IN_OBUF(m1_oper1_rdata_int[20]),.OUT_OBUF(m1_m1_oper_in[20]));

	OBUF QL_INST_F2A_B_22_9 (.IN_OBUF(m1_oper1_rdata_int[19]),.OUT_OBUF(m1_m1_oper_in[19]));

	OBUF QL_INST_F2A_B_22_10 (.IN_OBUF(m1_oper1_rdata_int[18]),.OUT_OBUF(m1_m1_oper_in[18]));

	OBUF QL_INST_F2A_B_22_11 (.IN_OBUF(m1_oper1_rdata_int[17]),.OUT_OBUF(m1_m1_oper_in[17]));

	OBUF QL_INST_F2A_B_22_12 (.IN_OBUF(m1_oper1_rdata_int[16]),.OUT_OBUF(m1_m1_oper_in[16]));

	OBUF QL_INST_F2A_B_22_13 (.IN_OBUF(m1_oper1_rdata_int[15]),.OUT_OBUF(m1_m1_oper_in[15]));

	OBUF QL_INST_F2A_B_22_14 (.IN_OBUF(m1_oper1_rdata_int[14]),.OUT_OBUF(m1_m1_oper_in[14]));

	OBUF QL_INST_F2A_B_22_15 (.IN_OBUF(m1_oper1_rdata_int[13]),.OUT_OBUF(m1_m1_oper_in[13]));

	OBUF QL_INST_F2A_B_22_16 (.IN_OBUF(m1_oper1_rdata_int[12]),.OUT_OBUF(m1_m1_oper_in[12]));

	OBUF QL_INST_F2A_B_22_17 (.IN_OBUF(m1_oper1_rdata_int[11]),.OUT_OBUF(m1_m1_oper_in[11]));

	IBUF QL_INST_A2F_B_22_0 (.IN_IBUF(m1_m1_dataout[10]),.OUT_IBUF(m1_m1_dataout_int[10]));

	IBUF QL_INST_A2F_B_22_1 (.IN_IBUF(m1_m1_dataout[9]),.OUT_IBUF(m1_m1_dataout_int[9]));

	IBUF QL_INST_A2F_B_22_2 (.IN_IBUF(m1_m1_dataout[8]),.OUT_IBUF(m1_m1_dataout_int[8]));

	IBUF QL_INST_A2F_B_22_3 (.IN_IBUF(m1_m1_dataout[7]),.OUT_IBUF(m1_m1_dataout_int[7]));

	IBUF QL_INST_A2F_B_22_4 (.IN_IBUF(m1_m1_dataout[6]),.OUT_IBUF(m1_m1_dataout_int[6]));

	IBUF QL_INST_A2F_B_22_5 (.IN_IBUF(m1_m1_dataout[5]),.OUT_IBUF(m1_m1_dataout_int[5]));

	OBUF QL_INST_F2A_B_23_0 (.IN_OBUF(m1_oper1_rdata_int[10]),.OUT_OBUF(m1_m1_oper_in[10]));

	OBUF QL_INST_F2A_B_23_1 (.IN_OBUF(m1_oper1_rdata_int[9]),.OUT_OBUF(m1_m1_oper_in[9]));

	OBUF QL_INST_F2A_B_23_2 (.IN_OBUF(m1_oper1_rdata_int[8]),.OUT_OBUF(m1_m1_oper_in[8]));

	OBUF QL_INST_F2A_B_23_3 (.IN_OBUF(m1_oper1_rdata_int[7]),.OUT_OBUF(m1_m1_oper_in[7]));

	OBUF QL_INST_F2A_B_23_4 (.IN_OBUF(m1_oper1_rdata_int[6]),.OUT_OBUF(m1_m1_oper_in[6]));

	OBUF QL_INST_F2A_B_23_5 (.IN_OBUF(m1_oper1_rdata_int[5]),.OUT_OBUF(m1_m1_oper_in[5]));

	OBUF QL_INST_F2A_B_23_6 (.IN_OBUF(m1_oper1_rdata_int[4]),.OUT_OBUF(m1_m1_oper_in[4]));

	OBUF QL_INST_F2A_B_23_7 (.IN_OBUF(m1_oper1_rdata_int[3]),.OUT_OBUF(m1_m1_oper_in[3]));

	OBUF QL_INST_F2A_B_23_8 (.IN_OBUF(m1_oper1_rdata_int[2]),.OUT_OBUF(m1_m1_oper_in[2]));

	OBUF QL_INST_F2A_B_23_9 (.IN_OBUF(m1_oper1_rdata_int[1]),.OUT_OBUF(m1_m1_oper_in[1]));

	OBUF QL_INST_F2A_B_23_10 (.IN_OBUF(m1_oper1_rdata_int[0]),.OUT_OBUF(m1_m1_oper_in[0]));

	IBUF QL_INST_A2F_B_23_0 (.IN_IBUF(m1_m1_dataout[4]),.OUT_IBUF(m1_m1_dataout_int[4]));

	IBUF QL_INST_A2F_B_23_1 (.IN_IBUF(m1_m1_dataout[3]),.OUT_IBUF(m1_m1_dataout_int[3]));

	IBUF QL_INST_A2F_B_23_2 (.IN_IBUF(m1_m1_dataout[2]),.OUT_IBUF(m1_m1_dataout_int[2]));

	IBUF QL_INST_A2F_B_23_3 (.IN_IBUF(m1_m1_dataout[1]),.OUT_IBUF(m1_m1_dataout_int[1]));

	IBUF QL_INST_A2F_B_23_4 (.IN_IBUF(m1_m1_dataout[0]),.OUT_IBUF(m1_m1_dataout_int[0]));

	OBUF QL_INST_F2A_B_24_16 (.IN_OBUF(m1_oper1_wdata_dup_0[31]),.OUT_OBUF(m1_oper1_wdata[31]));

	OBUF QL_INST_F2A_B_24_17 (.IN_OBUF(m1_oper1_wdata_dup_0[30]),.OUT_OBUF(m1_oper1_wdata[30]));

	DBUF QL_INST_F2Adef_B_24_1 (.IN_DBUF(GND),.OUT_DBUF(m1_oper1_powerdn));

	OBUF QL_INST_F2A_B_25_0 (.IN_OBUF(m1_oper1_wdata_dup_0[29]),.OUT_OBUF(m1_oper1_wdata[29]));

	OBUF QL_INST_F2A_B_25_1 (.IN_OBUF(m1_oper1_wdata_dup_0[28]),.OUT_OBUF(m1_oper1_wdata[28]));

	OBUF QL_INST_F2A_B_25_2 (.IN_OBUF(m1_oper1_wdata_dup_0[27]),.OUT_OBUF(m1_oper1_wdata[27]));

	OBUF QL_INST_F2A_B_25_3 (.IN_OBUF(m1_oper1_wdata_dup_0[26]),.OUT_OBUF(m1_oper1_wdata[26]));

	OBUF QL_INST_F2A_B_25_4 (.IN_OBUF(m1_oper1_wdata_dup_0[25]),.OUT_OBUF(m1_oper1_wdata[25]));

	OBUF QL_INST_F2A_B_25_5 (.IN_OBUF(m1_oper1_wdata_dup_0[24]),.OUT_OBUF(m1_oper1_wdata[24]));

	OBUF QL_INST_F2A_B_25_6 (.IN_OBUF(m1_oper1_wdata_dup_0[23]),.OUT_OBUF(m1_oper1_wdata[23]));

	OBUF QL_INST_F2A_B_25_7 (.IN_OBUF(m1_oper1_wdata_dup_0[22]),.OUT_OBUF(m1_oper1_wdata[22]));

	OBUF QL_INST_F2A_B_25_8 (.IN_OBUF(m1_oper1_wdata_dup_0[21]),.OUT_OBUF(m1_oper1_wdata[21]));

	OBUF QL_INST_F2A_B_25_9 (.IN_OBUF(m1_oper1_wdata_dup_0[20]),.OUT_OBUF(m1_oper1_wdata[20]));

	OBUF QL_INST_F2A_B_25_10 (.IN_OBUF(m1_oper1_wdata_dup_0[19]),.OUT_OBUF(m1_oper1_wdata[19]));

	OBUF QL_INST_F2A_B_25_11 (.IN_OBUF(m1_oper1_wdata_dup_0[18]),.OUT_OBUF(m1_oper1_wdata[18]));

	IBUF QL_INST_A2F_B_25_1 (.IN_IBUF(m1_oper1_rdata[31]),.OUT_IBUF(m1_oper1_rdata_int[31]));

	IBUF QL_INST_A2F_B_25_2 (.IN_IBUF(m1_oper1_rdata[30]),.OUT_IBUF(m1_oper1_rdata_int[30]));

	IBUF QL_INST_A2F_B_25_3 (.IN_IBUF(m1_oper1_rdata[29]),.OUT_IBUF(m1_oper1_rdata_int[29]));

	IBUF QL_INST_A2F_B_25_4 (.IN_IBUF(m1_oper1_rdata[28]),.OUT_IBUF(m1_oper1_rdata_int[28]));

	IBUF QL_INST_A2F_B_25_5 (.IN_IBUF(m1_oper1_rdata[27]),.OUT_IBUF(m1_oper1_rdata_int[27]));

	OBUF QL_INST_F2A_B_26_0 (.IN_OBUF(m1_oper1_wdata_dup_0[17]),.OUT_OBUF(m1_oper1_wdata[17]));

	OBUF QL_INST_F2A_B_26_1 (.IN_OBUF(m1_oper1_wdata_dup_0[16]),.OUT_OBUF(m1_oper1_wdata[16]));

	OBUF QL_INST_F2A_B_26_2 (.IN_OBUF(m1_oper1_wdata_dup_0[15]),.OUT_OBUF(m1_oper1_wdata[15]));

	OBUF QL_INST_F2A_B_26_3 (.IN_OBUF(m1_oper1_wdata_dup_0[14]),.OUT_OBUF(m1_oper1_wdata[14]));

	OBUF QL_INST_F2A_B_26_4 (.IN_OBUF(m1_oper1_wdata_dup_0[13]),.OUT_OBUF(m1_oper1_wdata[13]));

	OBUF QL_INST_F2A_B_26_5 (.IN_OBUF(m1_oper1_wdata_dup_0[12]),.OUT_OBUF(m1_oper1_wdata[12]));

	OBUF QL_INST_F2A_B_26_6 (.IN_OBUF(m1_oper1_wdata_dup_0[11]),.OUT_OBUF(m1_oper1_wdata[11]));

	OBUF QL_INST_F2A_B_26_7 (.IN_OBUF(m1_oper1_wdata_dup_0[10]),.OUT_OBUF(m1_oper1_wdata[10]));

	OBUF QL_INST_F2A_B_26_8 (.IN_OBUF(m1_oper1_wdata_dup_0[9]),.OUT_OBUF(m1_oper1_wdata[9]));

	OBUF QL_INST_F2A_B_26_9 (.IN_OBUF(m1_oper1_wdata_dup_0[8]),.OUT_OBUF(m1_oper1_wdata[8]));

	OBUF QL_INST_F2A_B_26_10 (.IN_OBUF(m1_oper1_wdata_dup_0[7]),.OUT_OBUF(m1_oper1_wdata[7]));

	OBUF QL_INST_F2A_B_26_11 (.IN_OBUF(m1_oper1_wdata_dup_0[6]),.OUT_OBUF(m1_oper1_wdata[6]));

	OBUF QL_INST_F2A_B_26_12 (.IN_OBUF(m1_oper1_wdata_dup_0[5]),.OUT_OBUF(m1_oper1_wdata[5]));

	OBUF QL_INST_F2A_B_26_13 (.IN_OBUF(m1_oper1_wdata_dup_0[4]),.OUT_OBUF(m1_oper1_wdata[4]));

	OBUF QL_INST_F2A_B_26_14 (.IN_OBUF(m1_oper1_wdata_dup_0[3]),.OUT_OBUF(m1_oper1_wdata[3]));

	OBUF QL_INST_F2A_B_26_15 (.IN_OBUF(m1_oper1_wdata_dup_0[2]),.OUT_OBUF(m1_oper1_wdata[2]));

	OBUF QL_INST_F2A_B_26_16 (.IN_OBUF(m1_oper1_wdata_dup_0[1]),.OUT_OBUF(m1_oper1_wdata[1]));

	OBUF QL_INST_F2A_B_26_17 (.IN_OBUF(m1_oper1_wdata_dup_0[0]),.OUT_OBUF(m1_oper1_wdata[0]));

	IBUF QL_INST_A2F_B_26_0 (.IN_IBUF(m1_oper1_rdata[26]),.OUT_IBUF(m1_oper1_rdata_int[26]));

	IBUF QL_INST_A2F_B_26_1 (.IN_IBUF(m1_oper1_rdata[25]),.OUT_IBUF(m1_oper1_rdata_int[25]));

	IBUF QL_INST_A2F_B_26_2 (.IN_IBUF(m1_oper1_rdata[24]),.OUT_IBUF(m1_oper1_rdata_int[24]));

	IBUF QL_INST_A2F_B_26_3 (.IN_IBUF(m1_oper1_rdata[23]),.OUT_IBUF(m1_oper1_rdata_int[23]));

	IBUF QL_INST_A2F_B_26_4 (.IN_IBUF(m1_oper1_rdata[22]),.OUT_IBUF(m1_oper1_rdata_int[22]));

	IBUF QL_INST_A2F_B_26_5 (.IN_IBUF(m1_oper1_rdata[21]),.OUT_IBUF(m1_oper1_rdata_int[21]));

	IBUF QL_INST_A2F_B_26_6 (.IN_IBUF(m1_oper1_rdata[20]),.OUT_IBUF(m1_oper1_rdata_int[20]));

	IBUF QL_INST_A2F_B_26_7 (.IN_IBUF(m1_oper1_rdata[19]),.OUT_IBUF(m1_oper1_rdata_int[19]));

	OBUF QL_INST_F2A_B_27_0 (.IN_OBUF(m1_oper1_waddr_dup_0[11]),.OUT_OBUF(m1_oper1_waddr[11]));

	OBUF QL_INST_F2A_B_27_1 (.IN_OBUF(m1_oper1_waddr_dup_0[10]),.OUT_OBUF(m1_oper1_waddr[10]));

	OBUF QL_INST_F2A_B_27_2 (.IN_OBUF(m1_oper1_waddr_dup_0[9]),.OUT_OBUF(m1_oper1_waddr[9]));

	OBUF QL_INST_F2A_B_27_3 (.IN_OBUF(m1_oper1_waddr_dup_0[8]),.OUT_OBUF(m1_oper1_waddr[8]));

	OBUF QL_INST_F2A_B_27_4 (.IN_OBUF(m1_oper1_waddr_dup_0[7]),.OUT_OBUF(m1_oper1_waddr[7]));

	OBUF QL_INST_F2A_B_27_5 (.IN_OBUF(m1_oper1_waddr_dup_0[6]),.OUT_OBUF(m1_oper1_waddr[6]));

	OBUF QL_INST_F2A_B_27_6 (.IN_OBUF(m1_oper1_waddr_dup_0[5]),.OUT_OBUF(m1_oper1_waddr[5]));

	OBUF QL_INST_F2A_B_27_7 (.IN_OBUF(m1_oper1_waddr_dup_0[4]),.OUT_OBUF(m1_oper1_waddr[4]));

	OBUF QL_INST_F2A_B_27_8 (.IN_OBUF(m1_oper1_waddr_dup_0[3]),.OUT_OBUF(m1_oper1_waddr[3]));

	OBUF QL_INST_F2A_B_27_9 (.IN_OBUF(m1_oper1_waddr_dup_0[2]),.OUT_OBUF(m1_oper1_waddr[2]));

	OBUF QL_INST_F2A_B_27_10 (.IN_OBUF(m1_oper1_waddr_dup_0[1]),.OUT_OBUF(m1_oper1_waddr[1]));

	OBUF QL_INST_F2A_B_27_11 (.IN_OBUF(m1_oper1_waddr_dup_0[0]),.OUT_OBUF(m1_oper1_waddr[0]));

	IBUF QL_INST_A2F_B_27_0 (.IN_IBUF(m1_oper1_rdata[18]),.OUT_IBUF(m1_oper1_rdata_int[18]));

	IBUF QL_INST_A2F_B_27_1 (.IN_IBUF(m1_oper1_rdata[17]),.OUT_IBUF(m1_oper1_rdata_int[17]));

	IBUF QL_INST_A2F_B_27_2 (.IN_IBUF(m1_oper1_rdata[16]),.OUT_IBUF(m1_oper1_rdata_int[16]));

	IBUF QL_INST_A2F_B_27_3 (.IN_IBUF(m1_oper1_rdata[15]),.OUT_IBUF(m1_oper1_rdata_int[15]));

	IBUF QL_INST_A2F_B_27_4 (.IN_IBUF(m1_oper1_rdata[14]),.OUT_IBUF(m1_oper1_rdata_int[14]));

	IBUF QL_INST_A2F_B_27_5 (.IN_IBUF(m1_oper1_rdata[13]),.OUT_IBUF(m1_oper1_rdata_int[13]));

	OBUF QL_INST_F2A_B_28_0 (.IN_OBUF(CLK_int_0__CAND0_BRSBR_28_padClk),.OUT_OBUF(m1_oper1_wclk));

	OBUF QL_INST_F2A_B_28_1 (.IN_OBUF(m0_oper1_wmode_dup_0[1]),.OUT_OBUF(m1_oper1_wmode[1]));

	OBUF QL_INST_F2A_B_28_2 (.IN_OBUF(m0_oper1_wmode_dup_0[0]),.OUT_OBUF(m1_oper1_wmode[0]));

	OBUF QL_INST_F2A_B_28_3 (.IN_OBUF(m0_oper1_wdsel_dup_0),.OUT_OBUF(m1_oper1_wdsel));

	OBUF QL_INST_F2A_B_28_4 (.IN_OBUF(m1_oper1_we_dup_0),.OUT_OBUF(m1_oper1_we));

	OBUF QL_INST_F2A_B_28_15 (.IN_OBUF(m0_oper1_rmode_dup_0[1]),.OUT_OBUF(m1_oper1_rmode[1]));

	OBUF QL_INST_F2A_B_28_16 (.IN_OBUF(m0_oper1_rmode_dup_0[0]),.OUT_OBUF(m1_oper1_rmode[0]));

	OBUF QL_INST_F2A_B_28_17 (.IN_OBUF(m1_oper1_raddr_dup_0[11]),.OUT_OBUF(m1_oper1_raddr[11]));

	IBUF QL_INST_A2F_B_28_1 (.IN_IBUF(m1_oper1_rdata[12]),.OUT_IBUF(m1_oper1_rdata_int[12]));

	IBUF QL_INST_A2F_B_28_2 (.IN_IBUF(m1_oper1_rdata[11]),.OUT_IBUF(m1_oper1_rdata_int[11]));

	IBUF QL_INST_A2F_B_28_3 (.IN_IBUF(m1_oper1_rdata[10]),.OUT_IBUF(m1_oper1_rdata_int[10]));

	IBUF QL_INST_A2F_B_28_4 (.IN_IBUF(m1_oper1_rdata[9]),.OUT_IBUF(m1_oper1_rdata_int[9]));

	IBUF QL_INST_A2F_B_28_5 (.IN_IBUF(m1_oper1_rdata[8]),.OUT_IBUF(m1_oper1_rdata_int[8]));

	IBUF QL_INST_A2F_B_28_6 (.IN_IBUF(m1_oper1_rdata[7]),.OUT_IBUF(m1_oper1_rdata_int[7]));

	IBUF QL_INST_A2F_B_28_7 (.IN_IBUF(m1_oper1_rdata[6]),.OUT_IBUF(m1_oper1_rdata_int[6]));

	OBUF QL_INST_F2A_B_29_0 (.IN_OBUF(CLK_int_0__CAND0_BRSBR_29_padClk),.OUT_OBUF(m1_oper1_rclk));

	OBUF QL_INST_F2A_B_29_1 (.IN_OBUF(m1_oper1_raddr_dup_0[10]),.OUT_OBUF(m1_oper1_raddr[10]));

	OBUF QL_INST_F2A_B_29_2 (.IN_OBUF(m1_oper1_raddr_dup_0[9]),.OUT_OBUF(m1_oper1_raddr[9]));

	OBUF QL_INST_F2A_B_29_3 (.IN_OBUF(m1_oper1_raddr_dup_0[8]),.OUT_OBUF(m1_oper1_raddr[8]));

	OBUF QL_INST_F2A_B_29_4 (.IN_OBUF(m1_oper1_raddr_dup_0[7]),.OUT_OBUF(m1_oper1_raddr[7]));

	OBUF QL_INST_F2A_B_29_5 (.IN_OBUF(m1_oper1_raddr_dup_0[6]),.OUT_OBUF(m1_oper1_raddr[6]));

	OBUF QL_INST_F2A_B_29_6 (.IN_OBUF(m1_oper1_raddr_dup_0[5]),.OUT_OBUF(m1_oper1_raddr[5]));

	OBUF QL_INST_F2A_B_29_7 (.IN_OBUF(m1_oper1_raddr_dup_0[4]),.OUT_OBUF(m1_oper1_raddr[4]));

	OBUF QL_INST_F2A_B_29_8 (.IN_OBUF(m1_oper1_raddr_dup_0[3]),.OUT_OBUF(m1_oper1_raddr[3]));

	OBUF QL_INST_F2A_B_29_9 (.IN_OBUF(m1_oper1_raddr_dup_0[2]),.OUT_OBUF(m1_oper1_raddr[2]));

	OBUF QL_INST_F2A_B_29_10 (.IN_OBUF(m1_oper1_raddr_dup_0[1]),.OUT_OBUF(m1_oper1_raddr[1]));

	OBUF QL_INST_F2A_B_29_11 (.IN_OBUF(m1_oper1_raddr_dup_0[0]),.OUT_OBUF(m1_oper1_raddr[0]));

	IBUF QL_INST_A2F_B_29_0 (.IN_IBUF(m1_oper1_rdata[5]),.OUT_IBUF(m1_oper1_rdata_int[5]));

	IBUF QL_INST_A2F_B_29_1 (.IN_IBUF(m1_oper1_rdata[4]),.OUT_IBUF(m1_oper1_rdata_int[4]));

	IBUF QL_INST_A2F_B_29_2 (.IN_IBUF(m1_oper1_rdata[3]),.OUT_IBUF(m1_oper1_rdata_int[3]));

	IBUF QL_INST_A2F_B_29_3 (.IN_IBUF(m1_oper1_rdata[2]),.OUT_IBUF(m1_oper1_rdata_int[2]));

	IBUF QL_INST_A2F_B_29_4 (.IN_IBUF(m1_oper1_rdata[1]),.OUT_IBUF(m1_oper1_rdata_int[1]));

	IBUF QL_INST_A2F_B_29_5 (.IN_IBUF(m1_oper1_rdata[0]),.OUT_IBUF(m1_oper1_rdata_int[0]));

	OBUF QL_INST_F2A_L_2_0 (.IN_OBUF(fpgaio_out_dup_0[0]),.OUT_OBUF(fpgaio_out[0]));

	OBUF QL_INST_F2A_L_2_1 (.IN_OBUF(fpgaio_oe_dup_0[0]),.OUT_OBUF(fpgaio_oe[0]));

	OBUF QL_INST_F2A_L_2_2 (.IN_OBUF(fpgaio_out_dup_0[1]),.OUT_OBUF(fpgaio_out[1]));

	OBUF QL_INST_F2A_L_2_3 (.IN_OBUF(fpgaio_oe_dup_0[1]),.OUT_OBUF(fpgaio_oe[1]));

	OBUF QL_INST_F2A_L_2_4 (.IN_OBUF(fpgaio_out_dup_0[2]),.OUT_OBUF(fpgaio_out[2]));

	OBUF QL_INST_F2A_L_2_5 (.IN_OBUF(fpgaio_oe_dup_0[2]),.OUT_OBUF(fpgaio_oe[2]));

	OBUF QL_INST_F2A_L_2_6 (.IN_OBUF(fpgaio_out_dup_0[3]),.OUT_OBUF(fpgaio_out[3]));

	OBUF QL_INST_F2A_L_2_7 (.IN_OBUF(fpgaio_oe_dup_0[3]),.OUT_OBUF(fpgaio_oe[3]));

	OBUF QL_INST_F2A_L_2_8 (.IN_OBUF(fpgaio_in_int[0]),.OUT_OBUF(events_o[0]));

	DBUF QL_INST_F2Adef_L_2_0 (.IN_DBUF(VCC),.OUT_DBUF(version[0]));

	DBUF QL_INST_F2Adef_L_2_1 (.IN_DBUF(GND),.OUT_DBUF(version[1]));

	DBUF QL_INST_F2Adef_L_2_2 (.IN_DBUF(VCC),.OUT_DBUF(version[2]));

	DBUF QL_INST_F2Adef_L_2_3 (.IN_DBUF(GND),.OUT_DBUF(version[3]));

	DBUF QL_INST_F2Adef_L_2_4 (.IN_DBUF(VCC),.OUT_DBUF(version[4]));

	DBUF QL_INST_F2Adef_L_2_5 (.IN_DBUF(GND),.OUT_DBUF(version[5]));

	DBUF QL_INST_F2Adef_L_2_6 (.IN_DBUF(VCC),.OUT_DBUF(version[6]));

	IBUF QL_INST_A2F_L_2_0 (.IN_IBUF(fpgaio_in[0]),.OUT_IBUF(fpgaio_in_int[0]));

	IBUF QL_INST_A2F_L_2_1 (.IN_IBUF(fpgaio_in[1]),.OUT_IBUF(fpgaio_in_int[1]));

	IBUF QL_INST_A2F_L_2_2 (.IN_IBUF(fpgaio_in[2]),.OUT_IBUF(fpgaio_in_int[2]));

	IBUF QL_INST_A2F_L_2_3 (.IN_IBUF(fpgaio_in[3]),.OUT_IBUF(fpgaio_in_int[3]));

	IBUF QL_INST_A2F_L_2_4 (.IN_IBUF(RESET[3]),.OUT_IBUF(RESET_int[3]));

	OBUF QL_INST_F2A_L_3_0 (.IN_OBUF(fpgaio_out_dup_0[4]),.OUT_OBUF(fpgaio_out[4]));

	OBUF QL_INST_F2A_L_3_1 (.IN_OBUF(fpgaio_oe_dup_0[4]),.OUT_OBUF(fpgaio_oe[4]));

	OBUF QL_INST_F2A_L_3_2 (.IN_OBUF(fpgaio_out_dup_0[5]),.OUT_OBUF(fpgaio_out[5]));

	OBUF QL_INST_F2A_L_3_3 (.IN_OBUF(fpgaio_oe_dup_0[5]),.OUT_OBUF(fpgaio_oe[5]));

	OBUF QL_INST_F2A_L_3_4 (.IN_OBUF(fpgaio_out_dup_0[6]),.OUT_OBUF(fpgaio_out[6]));

	OBUF QL_INST_F2A_L_3_5 (.IN_OBUF(fpgaio_oe_dup_0[6]),.OUT_OBUF(fpgaio_oe[6]));

	OBUF QL_INST_F2A_L_3_6 (.IN_OBUF(fpgaio_out_dup_0[7]),.OUT_OBUF(fpgaio_out[7]));

	OBUF QL_INST_F2A_L_3_7 (.IN_OBUF(fpgaio_oe_dup_0[7]),.OUT_OBUF(fpgaio_oe[7]));

	OBUF QL_INST_F2A_L_3_8 (.IN_OBUF(fpgaio_in_int[1]),.OUT_OBUF(events_o[1]));

	IBUF QL_INST_A2F_L_3_0 (.IN_IBUF(fpgaio_in[4]),.OUT_IBUF(fpgaio_in_int[4]));

	IBUF QL_INST_A2F_L_3_1 (.IN_IBUF(fpgaio_in[5]),.OUT_IBUF(fpgaio_in_int[5]));

	IBUF QL_INST_A2F_L_3_2 (.IN_IBUF(fpgaio_in[6]),.OUT_IBUF(fpgaio_in_int[6]));

	IBUF QL_INST_A2F_L_3_3 (.IN_IBUF(fpgaio_in[7]),.OUT_IBUF(fpgaio_in_int[7]));

	IBUF QL_INST_A2F_L_3_4 (.IN_IBUF(fpgaio_in[8]),.OUT_IBUF(fpgaio_in_int[8]));

	IBUF QL_INST_A2F_L_3_5 (.IN_IBUF(fpgaio_in[9]),.OUT_IBUF(fpgaio_in_int[9]));

	OBUF QL_INST_F2A_L_4_0 (.IN_OBUF(fpgaio_out_dup_0[8]),.OUT_OBUF(fpgaio_out[8]));

	OBUF QL_INST_F2A_L_4_1 (.IN_OBUF(fpgaio_oe_dup_0[8]),.OUT_OBUF(fpgaio_oe[8]));

	OBUF QL_INST_F2A_L_4_2 (.IN_OBUF(fpgaio_out_dup_0[9]),.OUT_OBUF(fpgaio_out[9]));

	OBUF QL_INST_F2A_L_4_3 (.IN_OBUF(fpgaio_oe_dup_0[9]),.OUT_OBUF(fpgaio_oe[9]));

	OBUF QL_INST_F2A_L_4_4 (.IN_OBUF(fpgaio_out_dup_0[10]),.OUT_OBUF(fpgaio_out[10]));

	OBUF QL_INST_F2A_L_4_5 (.IN_OBUF(fpgaio_oe_dup_0[10]),.OUT_OBUF(fpgaio_oe[10]));

	OBUF QL_INST_F2A_L_4_6 (.IN_OBUF(fpgaio_out_dup_0[11]),.OUT_OBUF(fpgaio_out[11]));

	OBUF QL_INST_F2A_L_4_7 (.IN_OBUF(fpgaio_oe_dup_0[11]),.OUT_OBUF(fpgaio_oe[11]));

	OBUF QL_INST_F2A_L_4_8 (.IN_OBUF(fpgaio_in_int[2]),.OUT_OBUF(events_o[2]));

	OBUF QL_INST_F2A_L_4_9 (.IN_OBUF(fpgaio_out_dup_0[12]),.OUT_OBUF(fpgaio_out[12]));

	OBUF QL_INST_F2A_L_4_10 (.IN_OBUF(fpgaio_oe_dup_0[12]),.OUT_OBUF(fpgaio_oe[12]));

	OBUF QL_INST_F2A_L_4_11 (.IN_OBUF(fpgaio_out_dup_0[13]),.OUT_OBUF(fpgaio_out[13]));

	OBUF QL_INST_F2A_L_4_12 (.IN_OBUF(fpgaio_oe_dup_0[13]),.OUT_OBUF(fpgaio_oe[13]));

	OBUF QL_INST_F2A_L_4_13 (.IN_OBUF(fpgaio_out_dup_0[14]),.OUT_OBUF(fpgaio_out[14]));

	OBUF QL_INST_F2A_L_4_14 (.IN_OBUF(fpgaio_oe_dup_0[14]),.OUT_OBUF(fpgaio_oe[14]));

	DBUF QL_INST_F2Adef_L_4_0 (.IN_DBUF(GND),.OUT_DBUF(version[7]));

	IBUF QL_INST_A2F_L_4_2 (.IN_IBUF(fpgaio_in[10]),.OUT_IBUF(fpgaio_in_int[10]));

	IBUF QL_INST_A2F_L_4_3 (.IN_IBUF(fpgaio_in[11]),.OUT_IBUF(fpgaio_in_int[11]));

	IBUF QL_INST_A2F_L_4_4 (.IN_IBUF(fpgaio_in[12]),.OUT_IBUF(fpgaio_in_int[12]));

	IBUF QL_INST_A2F_L_4_5 (.IN_IBUF(fpgaio_in[13]),.OUT_IBUF(fpgaio_in_int[13]));

	IBUF QL_INST_A2F_L_4_6 (.IN_IBUF(fpgaio_in[14]),.OUT_IBUF(fpgaio_in_int[14]));

	IBUF QL_INST_A2F_L_4_7 (.IN_IBUF(fpgaio_in[15]),.OUT_IBUF(fpgaio_in_int[15]));

	OBUF QL_INST_F2A_L_5_0 (.IN_OBUF(fpgaio_out_dup_0[15]),.OUT_OBUF(fpgaio_out[15]));

	OBUF QL_INST_F2A_L_5_1 (.IN_OBUF(fpgaio_oe_dup_0[15]),.OUT_OBUF(fpgaio_oe[15]));

	OBUF QL_INST_F2A_L_5_2 (.IN_OBUF(fpgaio_in_int[3]),.OUT_OBUF(events_o[3]));

	OBUF QL_INST_F2A_L_5_3 (.IN_OBUF(fpgaio_out_dup_0[16]),.OUT_OBUF(fpgaio_out[16]));

	OBUF QL_INST_F2A_L_5_4 (.IN_OBUF(fpgaio_oe_dup_0[16]),.OUT_OBUF(fpgaio_oe[16]));

	OBUF QL_INST_F2A_L_5_5 (.IN_OBUF(fpgaio_out_dup_0[17]),.OUT_OBUF(fpgaio_out[17]));

	OBUF QL_INST_F2A_L_5_6 (.IN_OBUF(fpgaio_oe_dup_0[17]),.OUT_OBUF(fpgaio_oe[17]));

	OBUF QL_INST_F2A_L_5_7 (.IN_OBUF(fpgaio_out_dup_0[18]),.OUT_OBUF(fpgaio_out[18]));

	OBUF QL_INST_F2A_L_5_8 (.IN_OBUF(fpgaio_oe_dup_0[18]),.OUT_OBUF(fpgaio_oe[18]));

	OBUF QL_INST_F2A_L_5_9 (.IN_OBUF(fpgaio_out_dup_0[19]),.OUT_OBUF(fpgaio_out[19]));

	OBUF QL_INST_F2A_L_5_10 (.IN_OBUF(fpgaio_oe_dup_0[19]),.OUT_OBUF(fpgaio_oe[19]));

	OBUF QL_INST_F2A_L_5_11 (.IN_OBUF(fpgaio_in_int[4]),.OUT_OBUF(events_o[4]));

	IBUF QL_INST_A2F_L_5_0 (.IN_IBUF(fpgaio_in[16]),.OUT_IBUF(fpgaio_in_int[16]));

	IBUF QL_INST_A2F_L_5_1 (.IN_IBUF(fpgaio_in[17]),.OUT_IBUF(fpgaio_in_int[17]));

	IBUF QL_INST_A2F_L_5_2 (.IN_IBUF(fpgaio_in[18]),.OUT_IBUF(fpgaio_in_int[18]));

	IBUF QL_INST_A2F_L_5_3 (.IN_IBUF(fpgaio_in[19]),.OUT_IBUF(fpgaio_in_int[19]));

	IBUF QL_INST_A2F_L_5_4 (.IN_IBUF(fpgaio_in[20]),.OUT_IBUF(fpgaio_in_int[20]));

	IBUF QL_INST_A2F_L_5_5 (.IN_IBUF(fpgaio_in[21]),.OUT_IBUF(fpgaio_in_int[21]));

	OBUF QL_INST_F2A_L_6_0 (.IN_OBUF(fpgaio_out_dup_0[20]),.OUT_OBUF(fpgaio_out[20]));

	OBUF QL_INST_F2A_L_6_1 (.IN_OBUF(fpgaio_oe_dup_0[20]),.OUT_OBUF(fpgaio_oe[20]));

	OBUF QL_INST_F2A_L_6_2 (.IN_OBUF(fpgaio_out_dup_0[21]),.OUT_OBUF(fpgaio_out[21]));

	OBUF QL_INST_F2A_L_6_3 (.IN_OBUF(fpgaio_oe_dup_0[21]),.OUT_OBUF(fpgaio_oe[21]));

	OBUF QL_INST_F2A_L_6_4 (.IN_OBUF(fpgaio_out_dup_0[22]),.OUT_OBUF(fpgaio_out[22]));

	OBUF QL_INST_F2A_L_6_5 (.IN_OBUF(fpgaio_oe_dup_0[22]),.OUT_OBUF(fpgaio_oe[22]));

	OBUF QL_INST_F2A_L_6_6 (.IN_OBUF(fpgaio_out_dup_0[23]),.OUT_OBUF(fpgaio_out[23]));

	OBUF QL_INST_F2A_L_6_7 (.IN_OBUF(fpgaio_oe_dup_0[23]),.OUT_OBUF(fpgaio_oe[23]));

	OBUF QL_INST_F2A_L_6_8 (.IN_OBUF(fpgaio_in_int[5]),.OUT_OBUF(events_o[5]));

	OBUF QL_INST_F2A_L_6_9 (.IN_OBUF(fpgaio_out_dup_0[24]),.OUT_OBUF(fpgaio_out[24]));

	OBUF QL_INST_F2A_L_6_10 (.IN_OBUF(fpgaio_oe_dup_0[24]),.OUT_OBUF(fpgaio_oe[24]));

	OBUF QL_INST_F2A_L_6_11 (.IN_OBUF(fpgaio_out_dup_0[25]),.OUT_OBUF(fpgaio_out[25]));

	OBUF QL_INST_F2A_L_6_12 (.IN_OBUF(fpgaio_oe_dup_0[25]),.OUT_OBUF(fpgaio_oe[25]));

	OBUF QL_INST_F2A_L_6_13 (.IN_OBUF(fpgaio_out_dup_0[26]),.OUT_OBUF(fpgaio_out[26]));

	OBUF QL_INST_F2A_L_6_14 (.IN_OBUF(fpgaio_oe_dup_0[26]),.OUT_OBUF(fpgaio_oe[26]));

	OBUF QL_INST_F2A_L_6_15 (.IN_OBUF(fpgaio_out_dup_0[27]),.OUT_OBUF(fpgaio_out[27]));

	OBUF QL_INST_F2A_L_6_16 (.IN_OBUF(fpgaio_oe_dup_0[27]),.OUT_OBUF(fpgaio_oe[27]));

	OBUF QL_INST_F2A_L_6_17 (.IN_OBUF(fpgaio_in_int[6]),.OUT_OBUF(events_o[6]));

	IBUF QL_INST_A2F_L_6_0 (.IN_IBUF(fpgaio_in[22]),.OUT_IBUF(fpgaio_in_int[22]));

	IBUF QL_INST_A2F_L_6_1 (.IN_IBUF(fpgaio_in[23]),.OUT_IBUF(fpgaio_in_int[23]));

	IBUF QL_INST_A2F_L_6_2 (.IN_IBUF(fpgaio_in[24]),.OUT_IBUF(fpgaio_in_int[24]));

	IBUF QL_INST_A2F_L_6_3 (.IN_IBUF(fpgaio_in[25]),.OUT_IBUF(fpgaio_in_int[25]));

	IBUF QL_INST_A2F_L_6_4 (.IN_IBUF(fpgaio_in[26]),.OUT_IBUF(fpgaio_in_int[26]));

	IBUF QL_INST_A2F_L_6_5 (.IN_IBUF(fpgaio_in[27]),.OUT_IBUF(fpgaio_in_int[27]));

	IBUF QL_INST_A2F_L_7_0 (.IN_IBUF(fpgaio_in[28]),.OUT_IBUF(fpgaio_in_int[28]));

	IBUF QL_INST_A2F_L_7_1 (.IN_IBUF(fpgaio_in[29]),.OUT_IBUF(fpgaio_in_int[29]));

	IBUF QL_INST_A2F_L_7_2 (.IN_IBUF(fpgaio_in[30]),.OUT_IBUF(fpgaio_in_int[30]));

	IBUF QL_INST_A2F_L_7_3 (.IN_IBUF(fpgaio_in[31]),.OUT_IBUF(fpgaio_in_int[31]));

	IBUF QL_INST_A2F_L_7_4 (.IN_IBUF(lint_WDATA[0]),.OUT_IBUF(lint_WDATA_int[0]));

	IBUF QL_INST_A2F_L_7_5 (.IN_IBUF(lint_WDATA[1]),.OUT_IBUF(lint_WDATA_int[1]));

	OBUF QL_INST_F2A_L_8_0 (.IN_OBUF(fpgaio_out_dup_0[28]),.OUT_OBUF(fpgaio_out[28]));

	OBUF QL_INST_F2A_L_8_1 (.IN_OBUF(fpgaio_oe_dup_0[28]),.OUT_OBUF(fpgaio_oe[28]));

	OBUF QL_INST_F2A_L_8_2 (.IN_OBUF(fpgaio_out_dup_0[29]),.OUT_OBUF(fpgaio_out[29]));

	OBUF QL_INST_F2A_L_8_3 (.IN_OBUF(fpgaio_oe_dup_0[29]),.OUT_OBUF(fpgaio_oe[29]));

	OBUF QL_INST_F2A_L_8_4 (.IN_OBUF(fpgaio_out_dup_0[30]),.OUT_OBUF(fpgaio_out[30]));

	OBUF QL_INST_F2A_L_8_5 (.IN_OBUF(fpgaio_oe_dup_0[30]),.OUT_OBUF(fpgaio_oe[30]));

	OBUF QL_INST_F2A_L_8_6 (.IN_OBUF(fpgaio_out_dup_0[31]),.OUT_OBUF(fpgaio_out[31]));

	OBUF QL_INST_F2A_L_8_7 (.IN_OBUF(fpgaio_oe_dup_0[31]),.OUT_OBUF(fpgaio_oe[31]));

	OBUF QL_INST_F2A_L_8_8 (.IN_OBUF(fpgaio_in_int[7]),.OUT_OBUF(events_o[7]));

	IBUF QL_INST_A2F_L_8_0 (.IN_IBUF(lint_WDATA[2]),.OUT_IBUF(lint_WDATA_int[2]));

	IBUF QL_INST_A2F_L_8_1 (.IN_IBUF(lint_WDATA[3]),.OUT_IBUF(lint_WDATA_int[3]));

	IBUF QL_INST_A2F_L_8_2 (.IN_IBUF(lint_WDATA[4]),.OUT_IBUF(lint_WDATA_int[4]));

	IBUF QL_INST_A2F_L_8_3 (.IN_IBUF(lint_WDATA[5]),.OUT_IBUF(lint_WDATA_int[5]));

	IBUF QL_INST_A2F_L_8_4 (.IN_IBUF(lint_WDATA[6]),.OUT_IBUF(lint_WDATA_int[6]));

	IBUF QL_INST_A2F_L_8_5 (.IN_IBUF(lint_WDATA[7]),.OUT_IBUF(lint_WDATA_int[7]));

	IBUF QL_INST_A2F_L_8_6 (.IN_IBUF(lint_WDATA[8]),.OUT_IBUF(lint_WDATA_int[8]));

	IBUF QL_INST_A2F_L_8_7 (.IN_IBUF(lint_WDATA[9]),.OUT_IBUF(lint_WDATA_int[9]));

	IBUF QL_INST_A2F_L_9_0 (.IN_IBUF(lint_WDATA[10]),.OUT_IBUF(lint_WDATA_int[10]));

	IBUF QL_INST_A2F_L_9_1 (.IN_IBUF(lint_WDATA[11]),.OUT_IBUF(lint_WDATA_int[11]));

	IBUF QL_INST_A2F_L_9_2 (.IN_IBUF(lint_WDATA[12]),.OUT_IBUF(lint_WDATA_int[12]));

	IBUF QL_INST_A2F_L_9_3 (.IN_IBUF(lint_WDATA[13]),.OUT_IBUF(lint_WDATA_int[13]));

	IBUF QL_INST_A2F_L_9_4 (.IN_IBUF(lint_WDATA[14]),.OUT_IBUF(lint_WDATA_int[14]));

	IBUF QL_INST_A2F_L_9_5 (.IN_IBUF(lint_WDATA[15]),.OUT_IBUF(lint_WDATA_int[15]));

	IBUF QL_INST_A2F_L_10_0 (.IN_IBUF(lint_WDATA[16]),.OUT_IBUF(lint_WDATA_int[16]));

	IBUF QL_INST_A2F_L_10_1 (.IN_IBUF(lint_WDATA[17]),.OUT_IBUF(lint_WDATA_int[17]));

	IBUF QL_INST_A2F_L_10_2 (.IN_IBUF(lint_WDATA[18]),.OUT_IBUF(lint_WDATA_int[18]));

	IBUF QL_INST_A2F_L_10_3 (.IN_IBUF(lint_WDATA[19]),.OUT_IBUF(lint_WDATA_int[19]));

	IBUF QL_INST_A2F_L_10_4 (.IN_IBUF(lint_WDATA[20]),.OUT_IBUF(lint_WDATA_int[20]));

	IBUF QL_INST_A2F_L_10_5 (.IN_IBUF(lint_WDATA[21]),.OUT_IBUF(lint_WDATA_int[21]));

	IBUF QL_INST_A2F_L_10_6 (.IN_IBUF(lint_WDATA[22]),.OUT_IBUF(lint_WDATA_int[22]));

	IBUF QL_INST_A2F_L_10_7 (.IN_IBUF(lint_WDATA[23]),.OUT_IBUF(lint_WDATA_int[23]));

	IBUF QL_INST_A2F_L_11_0 (.IN_IBUF(lint_WDATA[24]),.OUT_IBUF(lint_WDATA_int[24]));

	IBUF QL_INST_A2F_L_11_1 (.IN_IBUF(lint_WDATA[25]),.OUT_IBUF(lint_WDATA_int[25]));

	IBUF QL_INST_A2F_L_11_2 (.IN_IBUF(lint_WDATA[26]),.OUT_IBUF(lint_WDATA_int[26]));

	IBUF QL_INST_A2F_L_11_3 (.IN_IBUF(lint_WDATA[27]),.OUT_IBUF(lint_WDATA_int[27]));

	IBUF QL_INST_A2F_L_11_4 (.IN_IBUF(lint_WDATA[28]),.OUT_IBUF(lint_WDATA_int[28]));

	IBUF QL_INST_A2F_L_11_5 (.IN_IBUF(lint_WDATA[29]),.OUT_IBUF(lint_WDATA_int[29]));

	OBUF QL_INST_F2A_L_12_8 (.IN_OBUF(lint_RDATA_dup_0[0]),.OUT_OBUF(lint_RDATA[0]));

	OBUF QL_INST_F2A_L_12_9 (.IN_OBUF(lint_RDATA_dup_0[1]),.OUT_OBUF(lint_RDATA[1]));

	OBUF QL_INST_F2A_L_12_10 (.IN_OBUF(lint_RDATA_dup_0[2]),.OUT_OBUF(lint_RDATA[2]));

	OBUF QL_INST_F2A_L_12_11 (.IN_OBUF(lint_RDATA_dup_0[3]),.OUT_OBUF(lint_RDATA[3]));

	OBUF QL_INST_F2A_L_12_12 (.IN_OBUF(lint_RDATA_dup_0[4]),.OUT_OBUF(lint_RDATA[4]));

	OBUF QL_INST_F2A_L_12_13 (.IN_OBUF(lint_RDATA_dup_0[5]),.OUT_OBUF(lint_RDATA[5]));

	OBUF QL_INST_F2A_L_12_14 (.IN_OBUF(lint_RDATA_dup_0[6]),.OUT_OBUF(lint_RDATA[6]));

	OBUF QL_INST_F2A_L_12_15 (.IN_OBUF(lint_RDATA_dup_0[7]),.OUT_OBUF(lint_RDATA[7]));

	OBUF QL_INST_F2A_L_12_16 (.IN_OBUF(lint_RDATA_dup_0[8]),.OUT_OBUF(lint_RDATA[8]));

	IBUF QL_INST_A2F_L_12_0 (.IN_IBUF(lint_WDATA[30]),.OUT_IBUF(lint_WDATA_int[30]));

	IBUF QL_INST_A2F_L_12_1 (.IN_IBUF(lint_WDATA[31]),.OUT_IBUF(lint_WDATA_int[31]));

	IBUF QL_INST_A2F_L_12_2 (.IN_IBUF(lint_REQ),.OUT_IBUF(lint_REQ_int));

	IBUF QL_INST_A2F_L_12_3 (.IN_IBUF(lint_WEN),.OUT_IBUF(lint_WEN_int));

	IBUF QL_INST_A2F_L_12_4 (.IN_IBUF(lint_BE[0]),.OUT_IBUF(lint_BE_int[0]));

	IBUF QL_INST_A2F_L_12_5 (.IN_IBUF(lint_BE[1]),.OUT_IBUF(lint_BE_int[1]));

	IBUF QL_INST_A2F_L_12_6 (.IN_IBUF(lint_BE[2]),.OUT_IBUF(lint_BE_int[2]));

	IBUF QL_INST_A2F_L_12_7 (.IN_IBUF(lint_BE[3]),.OUT_IBUF(lint_BE_int[3]));

	OBUF QL_INST_F2A_L_13_0 (.IN_OBUF(lint_RDATA_dup_0[9]),.OUT_OBUF(lint_RDATA[9]));

	OBUF QL_INST_F2A_L_13_1 (.IN_OBUF(lint_RDATA_dup_0[10]),.OUT_OBUF(lint_RDATA[10]));

	OBUF QL_INST_F2A_L_13_2 (.IN_OBUF(lint_RDATA_dup_0[11]),.OUT_OBUF(lint_RDATA[11]));

	OBUF QL_INST_F2A_L_13_3 (.IN_OBUF(lint_RDATA_dup_0[12]),.OUT_OBUF(lint_RDATA[12]));

	OBUF QL_INST_F2A_L_13_4 (.IN_OBUF(lint_RDATA_dup_0[13]),.OUT_OBUF(lint_RDATA[13]));

	OBUF QL_INST_F2A_L_13_5 (.IN_OBUF(lint_RDATA_dup_0[14]),.OUT_OBUF(lint_RDATA[14]));

	OBUF QL_INST_F2A_L_13_6 (.IN_OBUF(lint_RDATA_dup_0[15]),.OUT_OBUF(lint_RDATA[15]));

	IBUF QL_INST_A2F_L_13_0 (.IN_IBUF(lint_ADDR[0]),.OUT_IBUF(lint_ADDR_int[0]));

	IBUF QL_INST_A2F_L_13_1 (.IN_IBUF(lint_ADDR[1]),.OUT_IBUF(lint_ADDR_int[1]));

	IBUF QL_INST_A2F_L_13_2 (.IN_IBUF(lint_ADDR[2]),.OUT_IBUF(lint_ADDR_int[2]));

	IBUF QL_INST_A2F_L_13_3 (.IN_IBUF(lint_ADDR[3]),.OUT_IBUF(lint_ADDR_int[3]));

	IBUF QL_INST_A2F_L_13_4 (.IN_IBUF(lint_ADDR[4]),.OUT_IBUF(lint_ADDR_int[4]));

	IBUF QL_INST_A2F_L_13_5 (.IN_IBUF(lint_ADDR[5]),.OUT_IBUF(lint_ADDR_int[5]));

	OBUF QL_INST_F2A_L_14_0 (.IN_OBUF(CLK_int_0__CAND0_TLSBL_0_padClk),.OUT_OBUF(lint_clk));

	OBUF QL_INST_F2A_L_14_1 (.IN_OBUF(lint_RDATA_dup_0[16]),.OUT_OBUF(lint_RDATA[16]));

	OBUF QL_INST_F2A_L_14_2 (.IN_OBUF(lint_RDATA_dup_0[17]),.OUT_OBUF(lint_RDATA[17]));

	OBUF QL_INST_F2A_L_14_3 (.IN_OBUF(lint_RDATA_dup_0[18]),.OUT_OBUF(lint_RDATA[18]));

	OBUF QL_INST_F2A_L_14_4 (.IN_OBUF(lint_RDATA_dup_0[19]),.OUT_OBUF(lint_RDATA[19]));

	OBUF QL_INST_F2A_L_14_5 (.IN_OBUF(lint_RDATA_dup_0[20]),.OUT_OBUF(lint_RDATA[20]));

	OBUF QL_INST_F2A_L_14_6 (.IN_OBUF(lint_RDATA_dup_0[21]),.OUT_OBUF(lint_RDATA[21]));

	OBUF QL_INST_F2A_L_14_7 (.IN_OBUF(lint_RDATA_dup_0[22]),.OUT_OBUF(lint_RDATA[22]));

	OBUF QL_INST_F2A_L_14_8 (.IN_OBUF(lint_RDATA_dup_0[23]),.OUT_OBUF(lint_RDATA[23]));

	OBUF QL_INST_F2A_L_14_9 (.IN_OBUF(lint_VALID_dup_0),.OUT_OBUF(lint_VALID));

	IBUF QL_INST_A2F_L_14_0 (.IN_IBUF(lint_ADDR[6]),.OUT_IBUF(lint_ADDR_int[6]));

	IBUF QL_INST_A2F_L_14_1 (.IN_IBUF(lint_ADDR[7]),.OUT_IBUF(lint_ADDR_int[7]));

	IBUF QL_INST_A2F_L_14_2 (.IN_IBUF(lint_ADDR[8]),.OUT_IBUF(lint_ADDR_int[8]));

	IBUF QL_INST_A2F_L_14_3 (.IN_IBUF(lint_ADDR[9]),.OUT_IBUF(lint_ADDR_int[9]));

	IBUF QL_INST_A2F_L_14_4 (.IN_IBUF(lint_ADDR[10]),.OUT_IBUF(lint_ADDR_int[10]));

	IBUF QL_INST_A2F_L_14_5 (.IN_IBUF(lint_ADDR[11]),.OUT_IBUF(lint_ADDR_int[11]));

	IBUF QL_INST_A2F_L_14_6 (.IN_IBUF(lint_ADDR[12]),.OUT_IBUF(lint_ADDR_int[12]));

	IBUF QL_INST_A2F_L_14_7 (.IN_IBUF(lint_ADDR[13]),.OUT_IBUF(lint_ADDR_int[13]));

	OBUF QL_INST_F2A_L_15_0 (.IN_OBUF(lint_RDATA_dup_0[24]),.OUT_OBUF(lint_RDATA[24]));

	OBUF QL_INST_F2A_L_15_1 (.IN_OBUF(lint_RDATA_dup_0[25]),.OUT_OBUF(lint_RDATA[25]));

	OBUF QL_INST_F2A_L_15_2 (.IN_OBUF(lint_RDATA_dup_0[26]),.OUT_OBUF(lint_RDATA[26]));

	OBUF QL_INST_F2A_L_15_3 (.IN_OBUF(lint_RDATA_dup_0[27]),.OUT_OBUF(lint_RDATA[27]));

	OBUF QL_INST_F2A_L_15_4 (.IN_OBUF(lint_RDATA_dup_0[28]),.OUT_OBUF(lint_RDATA[28]));

	OBUF QL_INST_F2A_L_15_5 (.IN_OBUF(lint_RDATA_dup_0[29]),.OUT_OBUF(lint_RDATA[29]));

	OBUF QL_INST_F2A_L_15_6 (.IN_OBUF(lint_RDATA_dup_0[30]),.OUT_OBUF(lint_RDATA[30]));

	OBUF QL_INST_F2A_L_15_7 (.IN_OBUF(lint_RDATA_dup_0[31]),.OUT_OBUF(lint_RDATA[31]));

	OBUF QL_INST_F2A_L_15_8 (.IN_OBUF(lint_GNT_dup_0),.OUT_OBUF(lint_GNT));

	IBUF QL_INST_A2F_L_15_0 (.IN_IBUF(lint_ADDR[14]),.OUT_IBUF(lint_ADDR_int[14]));

	IBUF QL_INST_A2F_L_15_1 (.IN_IBUF(lint_ADDR[15]),.OUT_IBUF(lint_ADDR_int[15]));

	IBUF QL_INST_A2F_L_15_2 (.IN_IBUF(lint_ADDR[16]),.OUT_IBUF(lint_ADDR_int[16]));

	IBUF QL_INST_A2F_L_15_3 (.IN_IBUF(lint_ADDR[17]),.OUT_IBUF(lint_ADDR_int[17]));

	IBUF QL_INST_A2F_L_15_4 (.IN_IBUF(lint_ADDR[18]),.OUT_IBUF(lint_ADDR_int[18]));

	IBUF QL_INST_A2F_L_15_5 (.IN_IBUF(lint_ADDR[19]),.OUT_IBUF(lint_ADDR_int[19]));

	IBUF QL_INST_A2F_L_16_0 (.IN_IBUF(fpgaio_in[64]),.OUT_IBUF(fpgaio_in_int[64]));

	IBUF QL_INST_A2F_L_16_1 (.IN_IBUF(fpgaio_in[65]),.OUT_IBUF(fpgaio_in_int[65]));

	IBUF QL_INST_A2F_L_16_2 (.IN_IBUF(fpgaio_in[66]),.OUT_IBUF(fpgaio_in_int[66]));

	IBUF QL_INST_A2F_L_16_3 (.IN_IBUF(fpgaio_in[67]),.OUT_IBUF(fpgaio_in_int[67]));

	IBUF QL_INST_A2F_L_16_4 (.IN_IBUF(fpgaio_in[68]),.OUT_IBUF(fpgaio_in_int[68]));

	IBUF QL_INST_A2F_L_16_5 (.IN_IBUF(fpgaio_in[69]),.OUT_IBUF(fpgaio_in_int[69]));

	IBUF QL_INST_A2F_L_16_6 (.IN_IBUF(fpgaio_in[70]),.OUT_IBUF(fpgaio_in_int[70]));

	IBUF QL_INST_A2F_L_16_7 (.IN_IBUF(fpgaio_in[71]),.OUT_IBUF(fpgaio_in_int[71]));

	OBUF QL_INST_F2A_L_17_0 (.IN_OBUF(fpgaio_out_dup_0[64]),.OUT_OBUF(fpgaio_out[64]));

	OBUF QL_INST_F2A_L_17_1 (.IN_OBUF(fpgaio_oe_dup_0[64]),.OUT_OBUF(fpgaio_oe[64]));

	OBUF QL_INST_F2A_L_17_2 (.IN_OBUF(fpgaio_out_dup_0[65]),.OUT_OBUF(fpgaio_out[65]));

	OBUF QL_INST_F2A_L_17_3 (.IN_OBUF(fpgaio_oe_dup_0[65]),.OUT_OBUF(fpgaio_oe[65]));

	OBUF QL_INST_F2A_L_17_4 (.IN_OBUF(fpgaio_out_dup_0[66]),.OUT_OBUF(fpgaio_out[66]));

	OBUF QL_INST_F2A_L_17_5 (.IN_OBUF(fpgaio_oe_dup_0[66]),.OUT_OBUF(fpgaio_oe[66]));

	OBUF QL_INST_F2A_L_17_6 (.IN_OBUF(fpgaio_out_dup_0[67]),.OUT_OBUF(fpgaio_out[67]));

	OBUF QL_INST_F2A_L_17_7 (.IN_OBUF(fpgaio_oe_dup_0[67]),.OUT_OBUF(fpgaio_oe[67]));

	IBUF QL_INST_A2F_L_17_0 (.IN_IBUF(fpgaio_in[72]),.OUT_IBUF(fpgaio_in_int[72]));

	IBUF QL_INST_A2F_L_17_1 (.IN_IBUF(fpgaio_in[73]),.OUT_IBUF(fpgaio_in_int[73]));

	IBUF QL_INST_A2F_L_17_2 (.IN_IBUF(fpgaio_in[74]),.OUT_IBUF(fpgaio_in_int[74]));

	IBUF QL_INST_A2F_L_17_3 (.IN_IBUF(fpgaio_in[75]),.OUT_IBUF(fpgaio_in_int[75]));

	IBUF QL_INST_A2F_L_17_4 (.IN_IBUF(fpgaio_in[76]),.OUT_IBUF(fpgaio_in_int[76]));

	IBUF QL_INST_A2F_L_17_5 (.IN_IBUF(fpgaio_in[77]),.OUT_IBUF(fpgaio_in_int[77]));

	OBUF QL_INST_F2A_L_18_0 (.IN_OBUF(fpgaio_out_dup_0[68]),.OUT_OBUF(fpgaio_out[68]));

	OBUF QL_INST_F2A_L_18_1 (.IN_OBUF(fpgaio_oe_dup_0[68]),.OUT_OBUF(fpgaio_oe[68]));

	OBUF QL_INST_F2A_L_18_2 (.IN_OBUF(fpgaio_out_dup_0[69]),.OUT_OBUF(fpgaio_out[69]));

	OBUF QL_INST_F2A_L_18_3 (.IN_OBUF(fpgaio_oe_dup_0[69]),.OUT_OBUF(fpgaio_oe[69]));

	OBUF QL_INST_F2A_L_18_4 (.IN_OBUF(fpgaio_out_dup_0[70]),.OUT_OBUF(fpgaio_out[70]));

	OBUF QL_INST_F2A_L_18_5 (.IN_OBUF(fpgaio_oe_dup_0[70]),.OUT_OBUF(fpgaio_oe[70]));

	OBUF QL_INST_F2A_L_18_6 (.IN_OBUF(fpgaio_out_dup_0[71]),.OUT_OBUF(fpgaio_out[71]));

	OBUF QL_INST_F2A_L_18_7 (.IN_OBUF(fpgaio_oe_dup_0[71]),.OUT_OBUF(fpgaio_oe[71]));

	OBUF QL_INST_F2A_L_18_8 (.IN_OBUF(fpgaio_out_dup_0[72]),.OUT_OBUF(fpgaio_out[72]));

	OBUF QL_INST_F2A_L_18_9 (.IN_OBUF(fpgaio_oe_dup_0[72]),.OUT_OBUF(fpgaio_oe[72]));

	OBUF QL_INST_F2A_L_18_10 (.IN_OBUF(fpgaio_out_dup_0[73]),.OUT_OBUF(fpgaio_out[73]));

	OBUF QL_INST_F2A_L_18_11 (.IN_OBUF(fpgaio_oe_dup_0[73]),.OUT_OBUF(fpgaio_oe[73]));

	OBUF QL_INST_F2A_L_18_12 (.IN_OBUF(fpgaio_out_dup_0[74]),.OUT_OBUF(fpgaio_out[74]));

	OBUF QL_INST_F2A_L_18_13 (.IN_OBUF(fpgaio_oe_dup_0[74]),.OUT_OBUF(fpgaio_oe[74]));

	OBUF QL_INST_F2A_L_18_14 (.IN_OBUF(fpgaio_out_dup_0[75]),.OUT_OBUF(fpgaio_out[75]));

	OBUF QL_INST_F2A_L_18_15 (.IN_OBUF(fpgaio_oe_dup_0[75]),.OUT_OBUF(fpgaio_oe[75]));

	IBUF QL_INST_A2F_L_18_0 (.IN_IBUF(fpgaio_in[78]),.OUT_IBUF(fpgaio_in_int[78]));

	IBUF QL_INST_A2F_L_18_1 (.IN_IBUF(fpgaio_in[79]),.OUT_IBUF(fpgaio_in_int[79]));

	OBUF QL_INST_F2A_L_19_0 (.IN_OBUF(fpgaio_out_dup_0[76]),.OUT_OBUF(fpgaio_out[76]));

	OBUF QL_INST_F2A_L_19_1 (.IN_OBUF(fpgaio_oe_dup_0[76]),.OUT_OBUF(fpgaio_oe[76]));

	OBUF QL_INST_F2A_L_19_2 (.IN_OBUF(fpgaio_out_dup_0[77]),.OUT_OBUF(fpgaio_out[77]));

	OBUF QL_INST_F2A_L_19_3 (.IN_OBUF(fpgaio_oe_dup_0[77]),.OUT_OBUF(fpgaio_oe[77]));

	OBUF QL_INST_F2A_L_19_4 (.IN_OBUF(fpgaio_out_dup_0[78]),.OUT_OBUF(fpgaio_out[78]));

	OBUF QL_INST_F2A_L_19_5 (.IN_OBUF(fpgaio_oe_dup_0[78]),.OUT_OBUF(fpgaio_oe[78]));

	OBUF QL_INST_F2A_L_19_6 (.IN_OBUF(fpgaio_out_dup_0[79]),.OUT_OBUF(fpgaio_out[79]));

	OBUF QL_INST_F2A_L_19_7 (.IN_OBUF(fpgaio_oe_dup_0[79]),.OUT_OBUF(fpgaio_oe[79]));

	IBUF QL_INST_A2F_L_19_0 (.IN_IBUF(control_in[0]),.OUT_IBUF(control_in_int[0]));

	IBUF QL_INST_A2F_L_19_1 (.IN_IBUF(control_in[1]),.OUT_IBUF(control_in_int[1]));

	IBUF QL_INST_A2F_L_19_2 (.IN_IBUF(control_in[2]),.OUT_IBUF(control_in_int[2]));

	IBUF QL_INST_A2F_L_19_3 (.IN_IBUF(control_in[3]),.OUT_IBUF(control_in_int[3]));

	IBUF QL_INST_A2F_L_19_4 (.IN_IBUF(control_in[4]),.OUT_IBUF(control_in_int[4]));

	IBUF QL_INST_A2F_L_19_5 (.IN_IBUF(control_in[5]),.OUT_IBUF(control_in_int[5]));

	OBUF QL_INST_F2A_L_20_0 (.IN_OBUF(status_out_dup_0[0]),.OUT_OBUF(status_out[0]));

	OBUF QL_INST_F2A_L_20_1 (.IN_OBUF(status_out_dup_0[1]),.OUT_OBUF(status_out[1]));

	OBUF QL_INST_F2A_L_20_2 (.IN_OBUF(status_out_dup_0[2]),.OUT_OBUF(status_out[2]));

	OBUF QL_INST_F2A_L_20_3 (.IN_OBUF(status_out_dup_0[3]),.OUT_OBUF(status_out[3]));

	OBUF QL_INST_F2A_L_20_4 (.IN_OBUF(status_out_dup_0[4]),.OUT_OBUF(status_out[4]));

	OBUF QL_INST_F2A_L_20_5 (.IN_OBUF(status_out_dup_0[5]),.OUT_OBUF(status_out[5]));

	OBUF QL_INST_F2A_L_20_6 (.IN_OBUF(status_out_dup_0[6]),.OUT_OBUF(status_out[6]));

	OBUF QL_INST_F2A_L_20_7 (.IN_OBUF(status_out_dup_0[7]),.OUT_OBUF(status_out[7]));

	OBUF QL_INST_F2A_L_20_8 (.IN_OBUF(status_out_dup_0[8]),.OUT_OBUF(status_out[8]));

	OBUF QL_INST_F2A_L_20_9 (.IN_OBUF(status_out_dup_0[9]),.OUT_OBUF(status_out[9]));

	OBUF QL_INST_F2A_L_20_10 (.IN_OBUF(status_out_dup_0[10]),.OUT_OBUF(status_out[10]));

	OBUF QL_INST_F2A_L_20_11 (.IN_OBUF(status_out_dup_0[11]),.OUT_OBUF(status_out[11]));

	OBUF QL_INST_F2A_L_20_12 (.IN_OBUF(status_out_dup_0[12]),.OUT_OBUF(status_out[12]));

	OBUF QL_INST_F2A_L_20_13 (.IN_OBUF(status_out_dup_0[13]),.OUT_OBUF(status_out[13]));

	OBUF QL_INST_F2A_L_20_14 (.IN_OBUF(status_out_dup_0[14]),.OUT_OBUF(status_out[14]));

	OBUF QL_INST_F2A_L_20_15 (.IN_OBUF(status_out_dup_0[15]),.OUT_OBUF(status_out[15]));

	OBUF QL_INST_F2A_L_20_16 (.IN_OBUF(status_out_dup_0[16]),.OUT_OBUF(status_out[16]));

	OBUF QL_INST_F2A_L_20_17 (.IN_OBUF(status_out_dup_0[17]),.OUT_OBUF(status_out[17]));

	IBUF QL_INST_A2F_L_20_0 (.IN_IBUF(control_in[6]),.OUT_IBUF(control_in_int[6]));

	IBUF QL_INST_A2F_L_20_1 (.IN_IBUF(control_in[7]),.OUT_IBUF(control_in_int[7]));

	IBUF QL_INST_A2F_L_20_2 (.IN_IBUF(control_in[8]),.OUT_IBUF(control_in_int[8]));

	IBUF QL_INST_A2F_L_20_3 (.IN_IBUF(control_in[9]),.OUT_IBUF(control_in_int[9]));

	IBUF QL_INST_A2F_L_20_4 (.IN_IBUF(control_in[10]),.OUT_IBUF(control_in_int[10]));

	IBUF QL_INST_A2F_L_20_5 (.IN_IBUF(control_in[11]),.OUT_IBUF(control_in_int[11]));

	IBUF QL_INST_A2F_L_20_6 (.IN_IBUF(control_in[12]),.OUT_IBUF(control_in_int[12]));

	IBUF QL_INST_A2F_L_20_7 (.IN_IBUF(control_in[13]),.OUT_IBUF(control_in_int[13]));

	OBUF QL_INST_F2A_L_21_0 (.IN_OBUF(status_out_dup_0[18]),.OUT_OBUF(status_out[18]));

	OBUF QL_INST_F2A_L_21_1 (.IN_OBUF(status_out_dup_0[19]),.OUT_OBUF(status_out[19]));

	OBUF QL_INST_F2A_L_21_2 (.IN_OBUF(status_out_dup_0[20]),.OUT_OBUF(status_out[20]));

	OBUF QL_INST_F2A_L_21_3 (.IN_OBUF(status_out_dup_0[21]),.OUT_OBUF(status_out[21]));

	OBUF QL_INST_F2A_L_21_4 (.IN_OBUF(status_out_dup_0[22]),.OUT_OBUF(status_out[22]));

	OBUF QL_INST_F2A_L_21_5 (.IN_OBUF(status_out_dup_0[23]),.OUT_OBUF(status_out[23]));

	OBUF QL_INST_F2A_L_21_6 (.IN_OBUF(status_out_dup_0[24]),.OUT_OBUF(status_out[24]));

	OBUF QL_INST_F2A_L_21_7 (.IN_OBUF(status_out_dup_0[25]),.OUT_OBUF(status_out[25]));

	OBUF QL_INST_F2A_L_21_8 (.IN_OBUF(status_out_dup_0[26]),.OUT_OBUF(status_out[26]));

	OBUF QL_INST_F2A_L_21_9 (.IN_OBUF(status_out_dup_0[27]),.OUT_OBUF(status_out[27]));

	OBUF QL_INST_F2A_L_21_10 (.IN_OBUF(status_out_dup_0[28]),.OUT_OBUF(status_out[28]));

	OBUF QL_INST_F2A_L_21_11 (.IN_OBUF(status_out_dup_0[29]),.OUT_OBUF(status_out[29]));

	IBUF QL_INST_A2F_L_21_0 (.IN_IBUF(control_in[14]),.OUT_IBUF(control_in_int[14]));

	IBUF QL_INST_A2F_L_21_1 (.IN_IBUF(control_in[15]),.OUT_IBUF(control_in_int[15]));

	IBUF QL_INST_A2F_L_21_2 (.IN_IBUF(control_in[16]),.OUT_IBUF(control_in_int[16]));

	IBUF QL_INST_A2F_L_21_3 (.IN_IBUF(control_in[17]),.OUT_IBUF(control_in_int[17]));

	IBUF QL_INST_A2F_L_21_4 (.IN_IBUF(control_in[18]),.OUT_IBUF(control_in_int[18]));

	IBUF QL_INST_A2F_L_21_5 (.IN_IBUF(control_in[19]),.OUT_IBUF(control_in_int[19]));

	OBUF QL_INST_F2A_L_22_0 (.IN_OBUF(status_out_dup_0[30]),.OUT_OBUF(status_out[30]));

	OBUF QL_INST_F2A_L_22_1 (.IN_OBUF(status_out_dup_0[31]),.OUT_OBUF(status_out[31]));

	IBUF QL_INST_A2F_L_22_0 (.IN_IBUF(control_in[20]),.OUT_IBUF(control_in_int[20]));

	IBUF QL_INST_A2F_L_22_1 (.IN_IBUF(control_in[21]),.OUT_IBUF(control_in_int[21]));

	IBUF QL_INST_A2F_L_22_2 (.IN_IBUF(control_in[22]),.OUT_IBUF(control_in_int[22]));

	IBUF QL_INST_A2F_L_22_3 (.IN_IBUF(control_in[23]),.OUT_IBUF(control_in_int[23]));

	IBUF QL_INST_A2F_L_22_4 (.IN_IBUF(control_in[24]),.OUT_IBUF(control_in_int[24]));

	IBUF QL_INST_A2F_L_22_5 (.IN_IBUF(control_in[25]),.OUT_IBUF(control_in_int[25]));

	IBUF QL_INST_A2F_L_22_6 (.IN_IBUF(control_in[26]),.OUT_IBUF(control_in_int[26]));

	IBUF QL_INST_A2F_L_23_0 (.IN_IBUF(control_in[27]),.OUT_IBUF(control_in_int[27]));

	IBUF QL_INST_A2F_L_23_1 (.IN_IBUF(control_in[28]),.OUT_IBUF(control_in_int[28]));

	IBUF QL_INST_A2F_L_23_2 (.IN_IBUF(control_in[29]),.OUT_IBUF(control_in_int[29]));

	IBUF QL_INST_A2F_L_23_3 (.IN_IBUF(control_in[30]),.OUT_IBUF(control_in_int[30]));

	IBUF QL_INST_A2F_L_23_4 (.IN_IBUF(control_in[31]),.OUT_IBUF(control_in_int[31]));

	OBUF QL_INST_F2A_L_25_0 (.IN_OBUF(fpgaio_out_dup_0[32]),.OUT_OBUF(fpgaio_out[32]));

	OBUF QL_INST_F2A_L_25_1 (.IN_OBUF(fpgaio_oe_dup_0[32]),.OUT_OBUF(fpgaio_oe[32]));

	OBUF QL_INST_F2A_L_25_2 (.IN_OBUF(fpgaio_out_dup_0[33]),.OUT_OBUF(fpgaio_out[33]));

	OBUF QL_INST_F2A_L_25_3 (.IN_OBUF(fpgaio_oe_dup_0[33]),.OUT_OBUF(fpgaio_oe[33]));

	OBUF QL_INST_F2A_L_25_4 (.IN_OBUF(fpgaio_out_dup_0[34]),.OUT_OBUF(fpgaio_out[34]));

	OBUF QL_INST_F2A_L_25_5 (.IN_OBUF(fpgaio_oe_dup_0[34]),.OUT_OBUF(fpgaio_oe[34]));

	OBUF QL_INST_F2A_L_25_6 (.IN_OBUF(fpgaio_out_dup_0[35]),.OUT_OBUF(fpgaio_out[35]));

	OBUF QL_INST_F2A_L_25_7 (.IN_OBUF(fpgaio_oe_dup_0[35]),.OUT_OBUF(fpgaio_oe[35]));

	OBUF QL_INST_F2A_L_25_8 (.IN_OBUF(fpgaio_in_int[8]),.OUT_OBUF(events_o[8]));

	IBUF QL_INST_A2F_L_25_0 (.IN_IBUF(fpgaio_in[32]),.OUT_IBUF(fpgaio_in_int[32]));

	IBUF QL_INST_A2F_L_25_1 (.IN_IBUF(fpgaio_in[33]),.OUT_IBUF(fpgaio_in_int[33]));

	IBUF QL_INST_A2F_L_25_2 (.IN_IBUF(RESET[2]),.OUT_IBUF(RESET_int[2]));

	IBUF QL_INST_A2F_L_25_3 (.IN_IBUF(fpgaio_in[34]),.OUT_IBUF(fpgaio_in_int[34]));

	IBUF QL_INST_A2F_L_25_4 (.IN_IBUF(fpgaio_in[35]),.OUT_IBUF(fpgaio_in_int[35]));

	OBUF QL_INST_F2A_L_26_0 (.IN_OBUF(fpgaio_out_dup_0[36]),.OUT_OBUF(fpgaio_out[36]));

	OBUF QL_INST_F2A_L_26_1 (.IN_OBUF(fpgaio_oe_dup_0[36]),.OUT_OBUF(fpgaio_oe[36]));

	OBUF QL_INST_F2A_L_26_2 (.IN_OBUF(fpgaio_out_dup_0[37]),.OUT_OBUF(fpgaio_out[37]));

	OBUF QL_INST_F2A_L_26_3 (.IN_OBUF(fpgaio_oe_dup_0[37]),.OUT_OBUF(fpgaio_oe[37]));

	OBUF QL_INST_F2A_L_26_4 (.IN_OBUF(fpgaio_out_dup_0[38]),.OUT_OBUF(fpgaio_out[38]));

	OBUF QL_INST_F2A_L_26_5 (.IN_OBUF(fpgaio_oe_dup_0[38]),.OUT_OBUF(fpgaio_oe[38]));

	OBUF QL_INST_F2A_L_26_6 (.IN_OBUF(fpgaio_out_dup_0[39]),.OUT_OBUF(fpgaio_out[39]));

	OBUF QL_INST_F2A_L_26_7 (.IN_OBUF(fpgaio_oe_dup_0[39]),.OUT_OBUF(fpgaio_oe[39]));

	OBUF QL_INST_F2A_L_26_8 (.IN_OBUF(fpgaio_in_int[9]),.OUT_OBUF(events_o[9]));

	IBUF QL_INST_A2F_L_26_0 (.IN_IBUF(fpgaio_in[36]),.OUT_IBUF(fpgaio_in_int[36]));

	IBUF QL_INST_A2F_L_26_1 (.IN_IBUF(fpgaio_in[37]),.OUT_IBUF(fpgaio_in_int[37]));

	IBUF QL_INST_A2F_L_26_2 (.IN_IBUF(fpgaio_in[38]),.OUT_IBUF(fpgaio_in_int[38]));

	IBUF QL_INST_A2F_L_26_3 (.IN_IBUF(fpgaio_in[39]),.OUT_IBUF(fpgaio_in_int[39]));

	OBUF QL_INST_F2A_L_27_0 (.IN_OBUF(fpgaio_out_dup_0[40]),.OUT_OBUF(fpgaio_out[40]));

	OBUF QL_INST_F2A_L_27_1 (.IN_OBUF(fpgaio_oe_dup_0[40]),.OUT_OBUF(fpgaio_oe[40]));

	OBUF QL_INST_F2A_L_27_2 (.IN_OBUF(fpgaio_out_dup_0[41]),.OUT_OBUF(fpgaio_out[41]));

	OBUF QL_INST_F2A_L_27_3 (.IN_OBUF(fpgaio_oe_dup_0[41]),.OUT_OBUF(fpgaio_oe[41]));

	OBUF QL_INST_F2A_L_27_4 (.IN_OBUF(fpgaio_out_dup_0[42]),.OUT_OBUF(fpgaio_out[42]));

	OBUF QL_INST_F2A_L_27_5 (.IN_OBUF(fpgaio_oe_dup_0[42]),.OUT_OBUF(fpgaio_oe[42]));

	OBUF QL_INST_F2A_L_27_6 (.IN_OBUF(fpgaio_out_dup_0[43]),.OUT_OBUF(fpgaio_out[43]));

	OBUF QL_INST_F2A_L_27_7 (.IN_OBUF(fpgaio_oe_dup_0[43]),.OUT_OBUF(fpgaio_oe[43]));

	OBUF QL_INST_F2A_L_27_8 (.IN_OBUF(fpgaio_in_int[10]),.OUT_OBUF(events_o[10]));

	IBUF QL_INST_A2F_L_27_0 (.IN_IBUF(fpgaio_in[40]),.OUT_IBUF(fpgaio_in_int[40]));

	IBUF QL_INST_A2F_L_27_1 (.IN_IBUF(fpgaio_in[41]),.OUT_IBUF(fpgaio_in_int[41]));

	IBUF QL_INST_A2F_L_27_2 (.IN_IBUF(fpgaio_in[42]),.OUT_IBUF(fpgaio_in_int[42]));

	IBUF QL_INST_A2F_L_27_3 (.IN_IBUF(fpgaio_in[43]),.OUT_IBUF(fpgaio_in_int[43]));

	OBUF QL_INST_F2A_L_28_0 (.IN_OBUF(fpgaio_out_dup_0[44]),.OUT_OBUF(fpgaio_out[44]));

	OBUF QL_INST_F2A_L_28_1 (.IN_OBUF(fpgaio_oe_dup_0[44]),.OUT_OBUF(fpgaio_oe[44]));

	OBUF QL_INST_F2A_L_28_2 (.IN_OBUF(fpgaio_out_dup_0[45]),.OUT_OBUF(fpgaio_out[45]));

	OBUF QL_INST_F2A_L_28_3 (.IN_OBUF(fpgaio_oe_dup_0[45]),.OUT_OBUF(fpgaio_oe[45]));

	OBUF QL_INST_F2A_L_28_4 (.IN_OBUF(fpgaio_out_dup_0[46]),.OUT_OBUF(fpgaio_out[46]));

	OBUF QL_INST_F2A_L_28_5 (.IN_OBUF(fpgaio_oe_dup_0[46]),.OUT_OBUF(fpgaio_oe[46]));

	OBUF QL_INST_F2A_L_28_6 (.IN_OBUF(fpgaio_out_dup_0[47]),.OUT_OBUF(fpgaio_out[47]));

	OBUF QL_INST_F2A_L_28_7 (.IN_OBUF(fpgaio_oe_dup_0[47]),.OUT_OBUF(fpgaio_oe[47]));

	OBUF QL_INST_F2A_L_28_8 (.IN_OBUF(fpgaio_in_int[11]),.OUT_OBUF(events_o[11]));

	IBUF QL_INST_A2F_L_28_0 (.IN_IBUF(fpgaio_in[44]),.OUT_IBUF(fpgaio_in_int[44]));

	IBUF QL_INST_A2F_L_28_1 (.IN_IBUF(fpgaio_in[45]),.OUT_IBUF(fpgaio_in_int[45]));

	IBUF QL_INST_A2F_L_28_2 (.IN_IBUF(fpgaio_in[46]),.OUT_IBUF(fpgaio_in_int[46]));

	IBUF QL_INST_A2F_L_28_3 (.IN_IBUF(fpgaio_in[47]),.OUT_IBUF(fpgaio_in_int[47]));

	OBUF QL_INST_F2A_L_29_0 (.IN_OBUF(fpgaio_out_dup_0[48]),.OUT_OBUF(fpgaio_out[48]));

	OBUF QL_INST_F2A_L_29_1 (.IN_OBUF(fpgaio_oe_dup_0[48]),.OUT_OBUF(fpgaio_oe[48]));

	OBUF QL_INST_F2A_L_29_2 (.IN_OBUF(fpgaio_out_dup_0[49]),.OUT_OBUF(fpgaio_out[49]));

	OBUF QL_INST_F2A_L_29_3 (.IN_OBUF(fpgaio_oe_dup_0[49]),.OUT_OBUF(fpgaio_oe[49]));

	OBUF QL_INST_F2A_L_29_4 (.IN_OBUF(fpgaio_out_dup_0[50]),.OUT_OBUF(fpgaio_out[50]));

	OBUF QL_INST_F2A_L_29_5 (.IN_OBUF(fpgaio_oe_dup_0[50]),.OUT_OBUF(fpgaio_oe[50]));

	OBUF QL_INST_F2A_L_29_6 (.IN_OBUF(fpgaio_out_dup_0[51]),.OUT_OBUF(fpgaio_out[51]));

	OBUF QL_INST_F2A_L_29_7 (.IN_OBUF(fpgaio_oe_dup_0[51]),.OUT_OBUF(fpgaio_oe[51]));

	OBUF QL_INST_F2A_L_29_8 (.IN_OBUF(fpgaio_in_int[12]),.OUT_OBUF(events_o[12]));

	IBUF QL_INST_A2F_L_29_0 (.IN_IBUF(fpgaio_in[48]),.OUT_IBUF(fpgaio_in_int[48]));

	IBUF QL_INST_A2F_L_29_1 (.IN_IBUF(fpgaio_in[49]),.OUT_IBUF(fpgaio_in_int[49]));

	IBUF QL_INST_A2F_L_29_2 (.IN_IBUF(fpgaio_in[50]),.OUT_IBUF(fpgaio_in_int[50]));

	IBUF QL_INST_A2F_L_29_3 (.IN_IBUF(fpgaio_in[51]),.OUT_IBUF(fpgaio_in_int[51]));

	OBUF QL_INST_F2A_L_30_0 (.IN_OBUF(fpgaio_out_dup_0[52]),.OUT_OBUF(fpgaio_out[52]));

	OBUF QL_INST_F2A_L_30_1 (.IN_OBUF(fpgaio_oe_dup_0[52]),.OUT_OBUF(fpgaio_oe[52]));

	OBUF QL_INST_F2A_L_30_2 (.IN_OBUF(fpgaio_out_dup_0[53]),.OUT_OBUF(fpgaio_out[53]));

	OBUF QL_INST_F2A_L_30_3 (.IN_OBUF(fpgaio_oe_dup_0[53]),.OUT_OBUF(fpgaio_oe[53]));

	OBUF QL_INST_F2A_L_30_4 (.IN_OBUF(fpgaio_out_dup_0[54]),.OUT_OBUF(fpgaio_out[54]));

	OBUF QL_INST_F2A_L_30_5 (.IN_OBUF(fpgaio_oe_dup_0[54]),.OUT_OBUF(fpgaio_oe[54]));

	OBUF QL_INST_F2A_L_30_6 (.IN_OBUF(fpgaio_out_dup_0[55]),.OUT_OBUF(fpgaio_out[55]));

	OBUF QL_INST_F2A_L_30_7 (.IN_OBUF(fpgaio_oe_dup_0[55]),.OUT_OBUF(fpgaio_oe[55]));

	OBUF QL_INST_F2A_L_30_8 (.IN_OBUF(fpgaio_in_int[13]),.OUT_OBUF(events_o[13]));

	IBUF QL_INST_A2F_L_30_0 (.IN_IBUF(fpgaio_in[52]),.OUT_IBUF(fpgaio_in_int[52]));

	IBUF QL_INST_A2F_L_30_1 (.IN_IBUF(fpgaio_in[53]),.OUT_IBUF(fpgaio_in_int[53]));

	IBUF QL_INST_A2F_L_30_2 (.IN_IBUF(fpgaio_in[54]),.OUT_IBUF(fpgaio_in_int[54]));

	IBUF QL_INST_A2F_L_30_3 (.IN_IBUF(fpgaio_in[55]),.OUT_IBUF(fpgaio_in_int[55]));

	OBUF QL_INST_F2A_L_31_0 (.IN_OBUF(fpgaio_out_dup_0[56]),.OUT_OBUF(fpgaio_out[56]));

	OBUF QL_INST_F2A_L_31_1 (.IN_OBUF(fpgaio_oe_dup_0[56]),.OUT_OBUF(fpgaio_oe[56]));

	OBUF QL_INST_F2A_L_31_2 (.IN_OBUF(fpgaio_out_dup_0[57]),.OUT_OBUF(fpgaio_out[57]));

	OBUF QL_INST_F2A_L_31_3 (.IN_OBUF(fpgaio_oe_dup_0[57]),.OUT_OBUF(fpgaio_oe[57]));

	OBUF QL_INST_F2A_L_31_4 (.IN_OBUF(fpgaio_out_dup_0[58]),.OUT_OBUF(fpgaio_out[58]));

	OBUF QL_INST_F2A_L_31_5 (.IN_OBUF(fpgaio_oe_dup_0[58]),.OUT_OBUF(fpgaio_oe[58]));

	OBUF QL_INST_F2A_L_31_6 (.IN_OBUF(fpgaio_out_dup_0[59]),.OUT_OBUF(fpgaio_out[59]));

	OBUF QL_INST_F2A_L_31_7 (.IN_OBUF(fpgaio_oe_dup_0[59]),.OUT_OBUF(fpgaio_oe[59]));

	OBUF QL_INST_F2A_L_31_8 (.IN_OBUF(fpgaio_in_int[14]),.OUT_OBUF(events_o[14]));

	IBUF QL_INST_A2F_L_31_0 (.IN_IBUF(fpgaio_in[56]),.OUT_IBUF(fpgaio_in_int[56]));

	IBUF QL_INST_A2F_L_31_1 (.IN_IBUF(fpgaio_in[57]),.OUT_IBUF(fpgaio_in_int[57]));

	IBUF QL_INST_A2F_L_31_2 (.IN_IBUF(fpgaio_in[58]),.OUT_IBUF(fpgaio_in_int[58]));

	IBUF QL_INST_A2F_L_31_3 (.IN_IBUF(fpgaio_in[59]),.OUT_IBUF(fpgaio_in_int[59]));

	OBUF QL_INST_F2A_L_32_0 (.IN_OBUF(fpgaio_out_dup_0[60]),.OUT_OBUF(fpgaio_out[60]));

	OBUF QL_INST_F2A_L_32_1 (.IN_OBUF(fpgaio_oe_dup_0[60]),.OUT_OBUF(fpgaio_oe[60]));

	OBUF QL_INST_F2A_L_32_2 (.IN_OBUF(fpgaio_out_dup_0[61]),.OUT_OBUF(fpgaio_out[61]));

	OBUF QL_INST_F2A_L_32_3 (.IN_OBUF(fpgaio_oe_dup_0[61]),.OUT_OBUF(fpgaio_oe[61]));

	OBUF QL_INST_F2A_L_32_4 (.IN_OBUF(fpgaio_out_dup_0[62]),.OUT_OBUF(fpgaio_out[62]));

	OBUF QL_INST_F2A_L_32_5 (.IN_OBUF(fpgaio_oe_dup_0[62]),.OUT_OBUF(fpgaio_oe[62]));

	OBUF QL_INST_F2A_L_32_6 (.IN_OBUF(fpgaio_out_dup_0[63]),.OUT_OBUF(fpgaio_out[63]));

	OBUF QL_INST_F2A_L_32_7 (.IN_OBUF(fpgaio_oe_dup_0[63]),.OUT_OBUF(fpgaio_oe[63]));

	OBUF QL_INST_F2A_L_32_8 (.IN_OBUF(fpgaio_in_int[15]),.OUT_OBUF(events_o[15]));

	IBUF QL_INST_A2F_L_32_0 (.IN_IBUF(fpgaio_in[60]),.OUT_IBUF(fpgaio_in_int[60]));

	IBUF QL_INST_A2F_L_32_1 (.IN_IBUF(fpgaio_in[61]),.OUT_IBUF(fpgaio_in_int[61]));

	IBUF QL_INST_A2F_L_32_2 (.IN_IBUF(fpgaio_in[62]),.OUT_IBUF(fpgaio_in_int[62]));

	IBUF QL_INST_A2F_L_32_3 (.IN_IBUF(fpgaio_in[63]),.OUT_IBUF(fpgaio_in_int[63]));

endmodule


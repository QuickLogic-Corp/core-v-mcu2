/*****************************************************************
          Vendor       : QuickLogic Corp.
          File Name    : top1.vq
          Author       : QuickLogic Corp.

          Description : Verilog Simulation Netlist file
******************************************************************/

`timescale 1ns / 10ps

module top1vq ( APB_CLK, CLK, RESET, events_o, fpgaio_in, fpgaio_oe, fpgaio_out, lint_ADDR, lint_BE, lint_GNT, lint_RDATA, lint_REQ, lint_VALID, lint_WDATA, lint_WEN, m0_coef_powerdn, m0_coef_raddr, m0_coef_rclk, m0_coef_rdata, m0_coef_rmode, m0_coef_waddr, m0_coef_wclk, m0_coef_wdata, m0_coef_wdsel, m0_coef_we, m0_coef_wmode, m0_m0_clk, m0_m0_clken, m0_m0_clr, m0_m0_coef_in, m0_m0_csel, m0_m0_dataout, m0_m0_mode, m0_m0_oper_in, m0_m0_osel, m0_m0_outsel, m0_m0_reset, m0_m0_rnd, m0_m0_sat, m0_m0_tc, m0_m1_clk, m0_m1_clken, m0_m1_clr, m0_m1_coef_in, m0_m1_csel, m0_m1_dataout, m0_m1_mode, m0_m1_oper_in, m0_m1_osel, m0_m1_outsel, m0_m1_reset, m0_m1_rnd, m0_m1_sat, m0_m1_tc, m0_oper0_powerdn, m0_oper0_raddr, m0_oper0_rclk, m0_oper0_rdata, m0_oper0_rmode, m0_oper0_waddr, m0_oper0_wclk, m0_oper0_wdata, m0_oper0_wdsel, m0_oper0_we, m0_oper0_wmode, m0_oper1_powerdn, m0_oper1_raddr, m0_oper1_rclk, m0_oper1_rdata, m0_oper1_rmode, m0_oper1_waddr, m0_oper1_wclk, m0_oper1_wdata, m0_oper1_wdsel, m0_oper1_we, m0_oper1_wmode, m1_coef_powerdn, m1_coef_raddr, m1_coef_rclk, m1_coef_rdata, m1_coef_rmode, m1_coef_waddr, m1_coef_wclk, m1_coef_wdata, m1_coef_wdsel, m1_coef_we, m1_coef_wmode, m1_m0_clk, m1_m0_clken, m1_m0_clr, m1_m0_coef_in, m1_m0_csel, m1_m0_dataout, m1_m0_mode, m1_m0_oper_in, m1_m0_osel, m1_m0_outsel, m1_m0_reset, m1_m0_rnd, m1_m0_sat, m1_m0_tc, m1_m1_clk, m1_m1_clken, m1_m1_clr, m1_m1_coef_in, m1_m1_csel, m1_m1_dataout, m1_m1_mode, m1_m1_oper_in, m1_m1_osel, m1_m1_outsel, m1_m1_reset, m1_m1_rnd, m1_m1_sat, m1_m1_tc, m1_oper0_powerdn, m1_oper0_raddr, m1_oper0_rclk, m1_oper0_rdata, m1_oper0_rmode, m1_oper0_waddr, m1_oper0_wclk, m1_oper0_wdata, m1_oper0_wdsel, m1_oper0_we, m1_oper0_wmode, m1_oper1_powerdn, m1_oper1_raddr, m1_oper1_rclk, m1_oper1_rdata, m1_oper1_rmode, m1_oper1_waddr, m1_oper1_wclk, m1_oper1_wdata, m1_oper1_wdsel, m1_oper1_we, m1_oper1_wmode, tcdm_addr_p0, tcdm_addr_p1, tcdm_addr_p2, tcdm_addr_p3, tcdm_be_p0, tcdm_be_p1, tcdm_be_p2, tcdm_be_p3, tcdm_clk_p0, tcdm_clk_p1, tcdm_clk_p2, tcdm_clk_p3, tcdm_gnt_p0, tcdm_gnt_p1, tcdm_gnt_p2, tcdm_gnt_p3, tcdm_rdata_p0, tcdm_rdata_p1, tcdm_rdata_p2, tcdm_rdata_p3, tcdm_req_p0, tcdm_req_p1, tcdm_req_p2, tcdm_req_p3, tcdm_valid_p0, tcdm_valid_p1, tcdm_valid_p2, tcdm_valid_p3, tcdm_wdata_p0, tcdm_wdata_p1, tcdm_wdata_p2, tcdm_wdata_p3, tcdm_we_p0, tcdm_we_p1, tcdm_we_p2, tcdm_we_p3);
output APB_CLK;
input [5:0] CLK;
input [3:0] RESET;
output [15:0] events_o;
input [79:0] fpgaio_in;
output [79:0] fpgaio_oe;
output [79:0] fpgaio_out;
input [19:0] lint_ADDR;
input [3:0] lint_BE;
output lint_GNT;
output [31:0] lint_RDATA;
input lint_REQ;
output lint_VALID;
input [31:0] lint_WDATA;
input lint_WEN;
output m0_coef_powerdn;
output [11:0] m0_coef_raddr;
output m0_coef_rclk;
input [31:0] m0_coef_rdata;
output [1:0] m0_coef_rmode;
output [11:0] m0_coef_waddr;
output m0_coef_wclk;
output [31:0] m0_coef_wdata;
output m0_coef_wdsel;
output m0_coef_we;
output [1:0] m0_coef_wmode;
output m0_m0_clk;
output m0_m0_clken;
output m0_m0_clr;
output [31:0] m0_m0_coef_in;
output m0_m0_csel;
input [31:0] m0_m0_dataout;
output [1:0] m0_m0_mode;
output [31:0] m0_m0_oper_in;
output m0_m0_osel;
output [5:0] m0_m0_outsel;
output m0_m0_reset;
output m0_m0_rnd;
output m0_m0_sat;
output m0_m0_tc;
output m0_m1_clk;
output m0_m1_clken;
output m0_m1_clr;
output [31:0] m0_m1_coef_in;
output m0_m1_csel;
input [31:0] m0_m1_dataout;
output [1:0] m0_m1_mode;
output [31:0] m0_m1_oper_in;
output m0_m1_osel;
output [5:0] m0_m1_outsel;
output m0_m1_reset;
output m0_m1_rnd;
output m0_m1_sat;
output m0_m1_tc;
output m0_oper0_powerdn;
output [11:0] m0_oper0_raddr;
output m0_oper0_rclk;
input [31:0] m0_oper0_rdata;
output [1:0] m0_oper0_rmode;
output [11:0] m0_oper0_waddr;
output m0_oper0_wclk;
output [31:0] m0_oper0_wdata;
output m0_oper0_wdsel;
output m0_oper0_we;
output [1:0] m0_oper0_wmode;
output m0_oper1_powerdn;
output [11:0] m0_oper1_raddr;
output m0_oper1_rclk;
input [31:0] m0_oper1_rdata;
output [1:0] m0_oper1_rmode;
output [11:0] m0_oper1_waddr;
output m0_oper1_wclk;
output [31:0] m0_oper1_wdata;
output m0_oper1_wdsel;
output m0_oper1_we;
output [1:0] m0_oper1_wmode;
output m1_coef_powerdn;
output [11:0] m1_coef_raddr;
output m1_coef_rclk;
input [31:0] m1_coef_rdata;
output [1:0] m1_coef_rmode;
output [11:0] m1_coef_waddr;
output m1_coef_wclk;
output [31:0] m1_coef_wdata;
output m1_coef_wdsel;
output m1_coef_we;
output [1:0] m1_coef_wmode;
output m1_m0_clk;
output m1_m0_clken;
output m1_m0_clr;
output [31:0] m1_m0_coef_in;
output m1_m0_csel;
input [31:0] m1_m0_dataout;
output [1:0] m1_m0_mode;
output [31:0] m1_m0_oper_in;
output m1_m0_osel;
output [5:0] m1_m0_outsel;
output m1_m0_reset;
output m1_m0_rnd;
output m1_m0_sat;
output m1_m0_tc;
output m1_m1_clk;
output m1_m1_clken;
output m1_m1_clr;
output [31:0] m1_m1_coef_in;
output m1_m1_csel;
input [31:0] m1_m1_dataout;
output [1:0] m1_m1_mode;
output [31:0] m1_m1_oper_in;
output m1_m1_osel;
output [5:0] m1_m1_outsel;
output m1_m1_reset;
output m1_m1_rnd;
output m1_m1_sat;
output m1_m1_tc;
output m1_oper0_powerdn;
output [11:0] m1_oper0_raddr;
output m1_oper0_rclk;
input [31:0] m1_oper0_rdata;
output [1:0] m1_oper0_rmode;
output [11:0] m1_oper0_waddr;
output m1_oper0_wclk;
output [31:0] m1_oper0_wdata;
output m1_oper0_wdsel;
output m1_oper0_we;
output [1:0] m1_oper0_wmode;
output m1_oper1_powerdn;
output [11:0] m1_oper1_raddr;
output m1_oper1_rclk;
input [31:0] m1_oper1_rdata;
output [1:0] m1_oper1_rmode;
output [11:0] m1_oper1_waddr;
output m1_oper1_wclk;
output [31:0] m1_oper1_wdata;
output m1_oper1_wdsel;
output m1_oper1_we;
output [1:0] m1_oper1_wmode;
output [19:0] tcdm_addr_p0;
output [19:0] tcdm_addr_p1;
output [19:0] tcdm_addr_p2;
output [19:0] tcdm_addr_p3;
output [3:0] tcdm_be_p0;
output [3:0] tcdm_be_p1;
output [3:0] tcdm_be_p2;
output [3:0] tcdm_be_p3;
output tcdm_clk_p0;
output tcdm_clk_p1;
output tcdm_clk_p2;
output tcdm_clk_p3;
input tcdm_gnt_p0;
input tcdm_gnt_p1;
input tcdm_gnt_p2;
input tcdm_gnt_p3;
input [31:0] tcdm_rdata_p0;
input [31:0] tcdm_rdata_p1;
input [31:0] tcdm_rdata_p2;
input [31:0] tcdm_rdata_p3;
output tcdm_req_p0;
output tcdm_req_p1;
output tcdm_req_p2;
output tcdm_req_p3;
input tcdm_valid_p0;
input tcdm_valid_p1;
input tcdm_valid_p2;
input tcdm_valid_p3;
output [31:0] tcdm_wdata_p0;
output [31:0] tcdm_wdata_p1;
output [31:0] tcdm_wdata_p2;
output [31:0] tcdm_wdata_p3;
output tcdm_we_p0;
output tcdm_we_p1;
output tcdm_we_p2;
output tcdm_we_p3;

supply1 VCC;
supply0 GND;

wire APB_CLK;
wire CLK_int_0__CAND0_BLSBL_1_padClk;
wire CLK_int_0__CAND0_BLSBL_2_padClk;
wire CLK_int_0__CAND0_BLSBL_3_padClk;
wire CLK_int_0__CAND0_BLSBL_4_padClk;
wire CLK_int_0__CAND0_BLSBL_5_padClk;
wire CLK_int_0__CAND0_BLSBL_6_padClk;
wire CLK_int_0__CAND0_BLSBL_7_padClk;
wire CLK_int_0__CAND0_BLSBL_8_padClk;
wire CLK_int_0__CAND0_BLSBR_10_padClk;
wire CLK_int_0__CAND0_BLSBR_11_padClk;
wire CLK_int_0__CAND0_BLSBR_13_padClk;
wire CLK_int_0__CAND0_BLSBR_14_padClk;
wire CLK_int_0__CAND0_BLSBR_15_padClk;
wire CLK_int_0__CAND0_BLSBR_16_padClk;
wire CLK_int_0__CAND0_BLSBR_9_padClk;
wire CLK_int_0__CAND0_BLSTL_0_padClk;
wire CLK_int_0__CAND0_BLSTL_1_padClk;
wire CLK_int_0__CAND0_BLSTL_3_padClk;
wire CLK_int_0__CAND0_BLSTL_4_padClk;
wire CLK_int_0__CAND0_BLSTL_5_padClk;
wire CLK_int_0__CAND0_BLSTL_6_padClk;
wire CLK_int_0__CAND0_BLSTL_7_padClk;
wire CLK_int_0__CAND0_BLSTL_8_padClk;
wire CLK_int_0__CAND0_BLSTR_10_padClk;
wire CLK_int_0__CAND0_BLSTR_11_padClk;
wire CLK_int_0__CAND0_BLSTR_12_padClk;
wire CLK_int_0__CAND0_BLSTR_13_padClk;
wire CLK_int_0__CAND0_BLSTR_14_padClk;
wire CLK_int_0__CAND0_BLSTR_15_padClk;
wire CLK_int_0__CAND0_BLSTR_16_padClk;
wire CLK_int_0__CAND0_BLSTR_9_padClk;
wire CLK_int_0__CAND0_BRSBL_17_padClk;
wire CLK_int_0__CAND0_BRSBL_18_padClk;
wire CLK_int_0__CAND0_BRSBL_19_padClk;
wire CLK_int_0__CAND0_BRSBL_23_padClk;
wire CLK_int_0__CAND0_BRSBL_24_padClk;
wire CLK_int_0__CAND0_BRSBR_25_padClk;
wire CLK_int_0__CAND0_BRSBR_26_padClk;
wire CLK_int_0__CAND0_BRSBR_27_padClk;
wire CLK_int_0__CAND0_BRSBR_28_padClk;
wire CLK_int_0__CAND0_BRSBR_29_padClk;
wire CLK_int_0__CAND0_BRSBR_30_padClk;
wire CLK_int_0__CAND0_BRSBR_31_padClk;
wire CLK_int_0__CAND0_BRSBR_32_padClk;
wire CLK_int_0__CAND0_BRSTL_17_padClk;
wire CLK_int_0__CAND0_BRSTL_18_padClk;
wire CLK_int_0__CAND0_BRSTL_19_padClk;
wire CLK_int_0__CAND0_BRSTL_20_padClk;
wire CLK_int_0__CAND0_BRSTL_21_padClk;
wire CLK_int_0__CAND0_BRSTL_22_padClk;
wire CLK_int_0__CAND0_BRSTR_28_padClk;
wire CLK_int_0__CAND0_BRSTR_29_padClk;
wire CLK_int_0__CAND0_BRSTR_30_padClk;
wire CLK_int_0__CAND0_BRSTR_31_padClk;
wire CLK_int_0__CAND0_BRSTR_32_padClk;
wire CLK_int_0__CAND0_BRSTR_33_padClk;
wire CLK_int_0__CAND0_TLSBL_1_padClk;
wire CLK_int_0__CAND0_TLSBL_3_padClk;
wire CLK_int_0__CAND0_TLSBL_4_padClk;
wire CLK_int_0__CAND0_TLSBL_5_padClk;
wire CLK_int_0__CAND0_TLSBL_6_padClk;
wire CLK_int_0__CAND0_TLSBL_7_padClk;
wire CLK_int_0__CAND0_TLSBL_8_padClk;
wire CLK_int_0__CAND0_TLSBR_10_padClk;
wire CLK_int_0__CAND0_TLSBR_11_padClk;
wire CLK_int_0__CAND0_TLSBR_12_padClk;
wire CLK_int_0__CAND0_TLSBR_13_padClk;
wire CLK_int_0__CAND0_TLSBR_14_padClk;
wire CLK_int_0__CAND0_TLSBR_15_padClk;
wire CLK_int_0__CAND0_TLSBR_16_padClk;
wire CLK_int_0__CAND0_TLSBR_9_padClk;
wire CLK_int_0__CAND0_TLSTL_1_padClk;
wire CLK_int_0__CAND0_TLSTL_2_padClk;
wire CLK_int_0__CAND0_TLSTL_3_padClk;
wire CLK_int_0__CAND0_TLSTL_4_padClk;
wire CLK_int_0__CAND0_TLSTL_5_padClk;
wire CLK_int_0__CAND0_TLSTL_6_padClk;
wire CLK_int_0__CAND0_TLSTL_7_padClk;
wire CLK_int_0__CAND0_TLSTL_8_padClk;
wire CLK_int_0__CAND0_TLSTR_12_padClk;
wire CLK_int_0__CAND0_TLSTR_13_padClk;
wire CLK_int_0__CAND0_TLSTR_14_padClk;
wire CLK_int_0__CAND0_TLSTR_15_padClk;
wire CLK_int_0__CAND0_TLSTR_16_padClk;
wire CLK_int_0__CAND0_TLSTR_9_padClk;
wire CLK_int_0__CAND0_TRSBL_17_padClk;
wire CLK_int_0__CAND0_TRSBL_18_padClk;
wire CLK_int_0__CAND0_TRSBL_19_padClk;
wire CLK_int_0__CAND0_TRSBL_20_padClk;
wire CLK_int_0__CAND0_TRSBL_21_padClk;
wire CLK_int_0__CAND0_TRSBL_22_padClk;
wire CLK_int_0__CAND0_TRSBR_29_padClk;
wire CLK_int_0__CAND0_TRSBR_30_padClk;
wire CLK_int_0__CAND0_TRSBR_31_padClk;
wire CLK_int_0__CAND0_TRSBR_32_padClk;
wire CLK_int_0__CAND0_TRSBR_33_padClk;
wire CLK_int_0__CAND0_TRSTL_17_padClk;
wire CLK_int_0__CAND0_TRSTL_18_padClk;
wire CLK_int_0__CAND0_TRSTL_19_padClk;
wire CLK_int_0__CAND0_TRSTL_23_padClk;
wire CLK_int_0__CAND0_TRSTL_24_padClk;
wire CLK_int_0__CAND0_TRSTR_25_padClk;
wire CLK_int_0__CAND0_TRSTR_26_padClk;
wire CLK_int_0__CAND0_TRSTR_27_padClk;
wire CLK_int_0__CAND0_TRSTR_28_padClk;
wire CLK_int_0__CAND0_TRSTR_29_padClk;
wire CLK_int_0__CAND0_TRSTR_30_padClk;
wire CLK_int_0__CAND0_TRSTR_31_padClk;
wire CLK_int_0__CAND0_TRSTR_32_padClk;
wire CLK_int_0__CAND0_TRSTR_33_padClk;
wire CLK_int_0__GMUX_0_padClk;
wire CLK_int_0__QMUX_BL0_padClk;
wire CLK_int_0__QMUX_BR0_padClk;
wire CLK_int_0__QMUX_TL0_padClk;
wire CLK_int_0__QMUX_TR0_padClk;
wire CLK_int_0__SQMUX_BLSBL0_padClk;
wire CLK_int_0__SQMUX_BLSBR0_padClk;
wire CLK_int_0__SQMUX_BLSTL0_padClk;
wire CLK_int_0__SQMUX_BLSTR0_padClk;
wire CLK_int_0__SQMUX_BRSBL0_padClk;
wire CLK_int_0__SQMUX_BRSBR0_padClk;
wire CLK_int_0__SQMUX_BRSTL0_padClk;
wire CLK_int_0__SQMUX_BRSTR0_padClk;
wire CLK_int_0__SQMUX_TLSBL0_padClk;
wire CLK_int_0__SQMUX_TLSBR0_padClk;
wire CLK_int_0__SQMUX_TLSTL0_padClk;
wire CLK_int_0__SQMUX_TLSTR0_padClk;
wire CLK_int_0__SQMUX_TRSBL0_padClk;
wire CLK_int_0__SQMUX_TRSBR0_padClk;
wire CLK_int_0__SQMUX_TRSTL0_padClk;
wire CLK_int_0__SQMUX_TRSTR0_padClk;
wire CLK_int_1__CAND1_TLSBL_8_padClk;
wire CLK_int_1__GMUX_1_padClk;
wire CLK_int_1__QMUX_TL1_padClk;
wire CLK_int_1__SQMUX_TLSBL1_padClk;
wire CLK_int_2__CAND2_TLSBL_8_padClk;
wire CLK_int_2__GMUX_2_padClk;
wire CLK_int_2__QMUX_TL2_padClk;
wire CLK_int_2__SQMUX_TLSBL2_padClk;
wire CLK_int_3__CAND3_BLSTL_6_padClk;
wire CLK_int_3__GMUX_3_padClk;
wire CLK_int_3__QMUX_BL3_padClk;
wire CLK_int_3__SQMUX_BLSTL3_padClk;
wire CLK_int_4__CAND4_TLSBL_8_padClk;
wire CLK_int_4__GMUX_4_padClk;
wire CLK_int_4__QMUX_TL4_padClk;
wire CLK_int_4__SQMUX_TLSBL4_padClk;
wire CLK_int_5__CAND5_TLSBL_7_padClk;
wire CLK_int_5__GMUX_5_padClk;
wire CLK_int_5__QMUX_TL5_padClk;
wire CLK_int_5__SQMUX_TLSBL5_padClk;
wire NET_0;
wire NET_1;
wire NET_10;
wire NET_100;
wire NET_101;
wire NET_102;
wire NET_103;
wire NET_104;
wire NET_105;
wire NET_106;
wire NET_107;
wire NET_108;
wire NET_109;
wire NET_11;
wire NET_110;
wire NET_110_CAND4_BRSTL_17_tpGCLKBUF;
wire NET_110_SQMUX_BRSTL4_tpGCLKBUF;
wire NET_111;
wire NET_112;
wire NET_113;
wire NET_114;
wire NET_115;
wire NET_116;
wire NET_117;
wire NET_118;
wire NET_119;
wire NET_12;
wire NET_120;
wire NET_121;
wire NET_122;
wire NET_123;
wire NET_124;
wire NET_124_CAND4_TLSBR_12_tpGCLKBUF;
wire NET_124_CAND4_TLSBR_13_tpGCLKBUF;
wire NET_124_CAND4_TLSBR_14_tpGCLKBUF;
wire NET_124_SQMUX_TLSBR4_tpGCLKBUF;
wire NET_125;
wire NET_125_CAND3_BRSTL_17_tpGCLKBUF;
wire NET_125_SQMUX_BRSTL3_tpGCLKBUF;
wire NET_126;
wire NET_127;
wire NET_128;
wire NET_129;
wire NET_13;
wire NET_130;
wire NET_131;
wire NET_132;
wire NET_133;
wire NET_134;
wire NET_135;
wire NET_136;
wire NET_137;
wire NET_138;
wire NET_139;
wire NET_14;
wire NET_140;
wire NET_141;
wire NET_142;
wire NET_143;
wire NET_144;
wire NET_145;
wire NET_146;
wire NET_147;
wire NET_148;
wire NET_149;
wire NET_15;
wire NET_150;
wire NET_151;
wire NET_152;
wire NET_153;
wire NET_154;
wire NET_155;
wire NET_156;
wire NET_157;
wire NET_158;
wire NET_159;
wire NET_15_CAND5_TLSBR_12_tpGCLKBUF;
wire NET_15_CAND5_TLSBR_13_tpGCLKBUF;
wire NET_15_CAND5_TLSBR_14_tpGCLKBUF;
wire NET_15_CAND5_TLSBR_15_tpGCLKBUF;
wire NET_15_CAND5_TLSBR_16_tpGCLKBUF;
wire NET_15_SQMUX_TLSBR5_tpGCLKBUF;
wire NET_16;
wire NET_160;
wire NET_161;
wire NET_162;
wire NET_163;
wire NET_164;
wire NET_165;
wire NET_166;
wire NET_167;
wire NET_168;
wire NET_169;
wire NET_17;
wire NET_170;
wire NET_171;
wire NET_172;
wire NET_173;
wire NET_174;
wire NET_175;
wire NET_176;
wire NET_177;
wire NET_178;
wire NET_179;
wire NET_17_CAND3_BLSTR_10_tpGCLKBUF;
wire NET_17_CAND3_BLSTR_11_tpGCLKBUF;
wire NET_17_CAND3_BLSTR_12_tpGCLKBUF;
wire NET_17_CAND3_BLSTR_13_tpGCLKBUF;
wire NET_17_CAND3_BLSTR_14_tpGCLKBUF;
wire NET_17_SQMUX_BLSTR3_tpGCLKBUF;
wire NET_18;
wire NET_180;
wire NET_181;
wire NET_182;
wire NET_183;
wire NET_184;
wire NET_185;
wire NET_186;
wire NET_187;
wire NET_188;
wire NET_189;
wire NET_18_CAND5_BLSTR_10_tpGCLKBUF;
wire NET_18_CAND5_BLSTR_11_tpGCLKBUF;
wire NET_18_CAND5_BLSTR_12_tpGCLKBUF;
wire NET_18_SQMUX_BLSTR5_tpGCLKBUF;
wire NET_19;
wire NET_190;
wire NET_191;
wire NET_192;
wire NET_193;
wire NET_194;
wire NET_195;
wire NET_196;
wire NET_197;
wire NET_198;
wire NET_199;
wire NET_2;
wire NET_20;
wire NET_200;
wire NET_201;
wire NET_202;
wire NET_203;
wire NET_204;
wire NET_205;
wire NET_206;
wire NET_207;
wire NET_208;
wire NET_209;
wire NET_21;
wire NET_210;
wire NET_211;
wire NET_212;
wire NET_213;
wire NET_214;
wire NET_215;
wire NET_216;
wire NET_217;
wire NET_218;
wire NET_219;
wire NET_22;
wire NET_220;
wire NET_221;
wire NET_222;
wire NET_223;
wire NET_224;
wire NET_225;
wire NET_226;
wire NET_227;
wire NET_228;
wire NET_229;
wire NET_23;
wire NET_230;
wire NET_231;
wire NET_232;
wire NET_233;
wire NET_234;
wire NET_235;
wire NET_236;
wire NET_237;
wire NET_238;
wire NET_239;
wire NET_24;
wire NET_240;
wire NET_241;
wire NET_242;
wire NET_243;
wire NET_244;
wire NET_245;
wire NET_246;
wire NET_247;
wire NET_248;
wire NET_249;
wire NET_25;
wire NET_250;
wire NET_251;
wire NET_252;
wire NET_253;
wire NET_254;
wire NET_255;
wire NET_256;
wire NET_257;
wire NET_258;
wire NET_259;
wire NET_26;
wire NET_260;
wire NET_261;
wire NET_262;
wire NET_263;
wire NET_264;
wire NET_265;
wire NET_266;
wire NET_267;
wire NET_268;
wire NET_269;
wire NET_27;
wire NET_270;
wire NET_271;
wire NET_272;
wire NET_273;
wire NET_274;
wire NET_275;
wire NET_276;
wire NET_277;
wire NET_278;
wire NET_279;
wire NET_28;
wire NET_280;
wire NET_281;
wire NET_282;
wire NET_283;
wire NET_284;
wire NET_285;
wire NET_286;
wire NET_287;
wire NET_288;
wire NET_289;
wire NET_28_CAND4_BLSTR_10_tpGCLKBUF;
wire NET_28_CAND4_BLSTR_11_tpGCLKBUF;
wire NET_28_CAND4_BLSTR_13_tpGCLKBUF;
wire NET_28_CAND4_BLSTR_14_tpGCLKBUF;
wire NET_28_CAND4_BLSTR_9_tpGCLKBUF;
wire NET_28_SQMUX_BLSTR4_tpGCLKBUF;
wire NET_29;
wire NET_290;
wire NET_291;
wire NET_292;
wire NET_293;
wire NET_294;
wire NET_295;
wire NET_296;
wire NET_297;
wire NET_298;
wire NET_299;
wire NET_29_CAND5_BLSTL_1_tpGCLKBUF;
wire NET_29_CAND5_BLSTL_7_tpGCLKBUF;
wire NET_29_CAND5_BLSTL_8_tpGCLKBUF;
wire NET_29_SQMUX_BLSTL5_tpGCLKBUF;
wire NET_3;
wire NET_30;
wire NET_300;
wire NET_301;
wire NET_302;
wire NET_303;
wire NET_304;
wire NET_305;
wire NET_306;
wire NET_307;
wire NET_308;
wire NET_309;
wire NET_31;
wire NET_310;
wire NET_311;
wire NET_312;
wire NET_313;
wire NET_314;
wire NET_315;
wire NET_316;
wire NET_317;
wire NET_318;
wire NET_319;
wire NET_32;
wire NET_320;
wire NET_321;
wire NET_322;
wire NET_323;
wire NET_324;
wire NET_325;
wire NET_326;
wire NET_327;
wire NET_328;
wire NET_329;
wire NET_32_CAND5_BLSBR_10_tpGCLKBUF;
wire NET_32_CAND5_BLSBR_11_tpGCLKBUF;
wire NET_32_CAND5_BLSBR_12_tpGCLKBUF;
wire NET_32_CAND5_BLSBR_13_tpGCLKBUF;
wire NET_32_SQMUX_BLSBR5_tpGCLKBUF;
wire NET_33;
wire NET_330;
wire NET_331;
wire NET_332;
wire NET_333;
wire NET_334;
wire NET_335;
wire NET_336;
wire NET_337;
wire NET_338;
wire NET_339;
wire NET_34;
wire NET_340;
wire NET_341;
wire NET_342;
wire NET_343;
wire NET_344;
wire NET_345;
wire NET_346;
wire NET_347;
wire NET_348;
wire NET_349;
wire NET_35;
wire NET_350;
wire NET_351;
wire NET_352;
wire NET_353;
wire NET_354;
wire NET_355;
wire NET_356;
wire NET_357;
wire NET_358;
wire NET_359;
wire NET_36;
wire NET_360;
wire NET_361;
wire NET_362;
wire NET_363;
wire NET_364;
wire NET_365;
wire NET_366;
wire NET_367;
wire NET_368;
wire NET_369;
wire NET_37;
wire NET_370;
wire NET_371;
wire NET_372;
wire NET_373;
wire NET_374;
wire NET_375;
wire NET_376;
wire NET_377;
wire NET_378;
wire NET_379;
wire NET_38;
wire NET_380;
wire NET_381;
wire NET_382;
wire NET_383;
wire NET_384;
wire NET_385;
wire NET_386;
wire NET_387;
wire NET_388;
wire NET_389;
wire NET_39;
wire NET_390;
wire NET_391;
wire NET_392;
wire NET_393;
wire NET_394;
wire NET_395;
wire NET_396;
wire NET_397;
wire NET_398;
wire NET_399;
wire NET_4;
wire NET_40;
wire NET_400;
wire NET_401;
wire NET_402;
wire NET_403;
wire NET_404;
wire NET_405;
wire NET_406;
wire NET_407;
wire NET_408;
wire NET_409;
wire NET_41;
wire NET_410;
wire NET_411;
wire NET_412;
wire NET_413;
wire NET_414;
wire NET_415;
wire NET_416;
wire NET_417;
wire NET_418;
wire NET_419;
wire NET_42;
wire NET_420;
wire NET_421;
wire NET_422;
wire NET_423;
wire NET_424;
wire NET_425;
wire NET_426;
wire NET_427;
wire NET_428;
wire NET_429;
wire NET_43;
wire NET_430;
wire NET_431;
wire NET_432;
wire NET_433;
wire NET_434;
wire NET_435;
wire NET_436;
wire NET_437;
wire NET_438;
wire NET_439;
wire NET_43_CAND3_BLSBR_11_tpGCLKBUF;
wire NET_43_CAND3_BLSBR_12_tpGCLKBUF;
wire NET_43_CAND3_BLSBR_13_tpGCLKBUF;
wire NET_43_CAND3_BLSBR_14_tpGCLKBUF;
wire NET_43_CAND3_BLSBR_15_tpGCLKBUF;
wire NET_43_SQMUX_BLSBR3_tpGCLKBUF;
wire NET_44;
wire NET_440;
wire NET_441;
wire NET_442;
wire NET_443;
wire NET_444;
wire NET_445;
wire NET_446;
wire NET_447;
wire NET_448;
wire NET_449;
wire NET_44_CAND4_BLSBR_12_tpGCLKBUF;
wire NET_44_CAND4_BLSBR_13_tpGCLKBUF;
wire NET_44_CAND4_BLSBR_14_tpGCLKBUF;
wire NET_44_CAND4_BLSBR_15_tpGCLKBUF;
wire NET_44_SQMUX_BLSBR4_tpGCLKBUF;
wire NET_45;
wire NET_450;
wire NET_451;
wire NET_452;
wire NET_453;
wire NET_454;
wire NET_455;
wire NET_456;
wire NET_457;
wire NET_458;
wire NET_459;
wire NET_46;
wire NET_460;
wire NET_461;
wire NET_462;
wire NET_463;
wire NET_464;
wire NET_465;
wire NET_466;
wire NET_467;
wire NET_468;
wire NET_469;
wire NET_46_CAND1_TLSTR_11_tpGCLKBUF;
wire NET_46_CAND1_TLSTR_12_tpGCLKBUF;
wire NET_46_CAND1_TLSTR_13_tpGCLKBUF;
wire NET_46_CAND1_TLSTR_14_tpGCLKBUF;
wire NET_46_CAND1_TLSTR_15_tpGCLKBUF;
wire NET_46_CAND1_TLSTR_16_tpGCLKBUF;
wire NET_46_SQMUX_TLSTR1_tpGCLKBUF;
wire NET_47;
wire NET_470;
wire NET_471;
wire NET_472;
wire NET_473;
wire NET_474;
wire NET_475;
wire NET_476;
wire NET_477;
wire NET_478;
wire NET_479;
wire NET_48;
wire NET_480;
wire NET_481;
wire NET_482;
wire NET_483;
wire NET_484;
wire NET_485;
wire NET_486;
wire NET_487;
wire NET_488;
wire NET_489;
wire NET_49;
wire NET_490;
wire NET_491;
wire NET_492;
wire NET_493;
wire NET_494;
wire NET_495;
wire NET_496;
wire NET_497;
wire NET_498;
wire NET_499;
wire NET_49_CAND4_TRSBL_17_tpGCLKBUF;
wire NET_49_CAND4_TRSBL_19_tpGCLKBUF;
wire NET_49_CAND4_TRSBL_20_tpGCLKBUF;
wire NET_49_CAND4_TRSBL_21_tpGCLKBUF;
wire NET_49_CAND4_TRSBL_22_tpGCLKBUF;
wire NET_49_SQMUX_TRSBL4_tpGCLKBUF;
wire NET_5;
wire NET_50;
wire NET_500;
wire NET_501;
wire NET_502;
wire NET_503;
wire NET_504;
wire NET_505;
wire NET_506;
wire NET_507;
wire NET_508;
wire NET_509;
wire NET_51;
wire NET_510;
wire NET_511;
wire NET_512;
wire NET_513;
wire NET_514;
wire NET_515;
wire NET_516;
wire NET_517;
wire NET_518;
wire NET_519;
wire NET_52;
wire NET_520;
wire NET_521;
wire NET_522;
wire NET_523;
wire NET_524;
wire NET_525;
wire NET_526;
wire NET_527;
wire NET_528;
wire NET_529;
wire NET_52_CAND2_TRSBL_18_tpGCLKBUF;
wire NET_52_CAND2_TRSBL_19_tpGCLKBUF;
wire NET_52_CAND2_TRSBL_20_tpGCLKBUF;
wire NET_52_CAND2_TRSBL_21_tpGCLKBUF;
wire NET_52_CAND2_TRSBL_22_tpGCLKBUF;
wire NET_52_SQMUX_TRSBL2_tpGCLKBUF;
wire NET_53;
wire NET_530;
wire NET_531;
wire NET_532;
wire NET_533;
wire NET_534;
wire NET_535;
wire NET_536;
wire NET_537;
wire NET_538;
wire NET_539;
wire NET_54;
wire NET_540;
wire NET_541;
wire NET_542;
wire NET_543;
wire NET_544;
wire NET_545;
wire NET_546;
wire NET_547;
wire NET_548;
wire NET_549;
wire NET_55;
wire NET_550;
wire NET_551;
wire NET_552;
wire NET_553;
wire NET_554;
wire NET_555;
wire NET_556;
wire NET_557;
wire NET_558;
wire NET_559;
wire NET_56;
wire NET_560;
wire NET_561;
wire NET_562;
wire NET_563;
wire NET_564;
wire NET_565;
wire NET_566;
wire NET_567;
wire NET_568;
wire NET_569;
wire NET_57;
wire NET_570;
wire NET_571;
wire NET_572;
wire NET_573;
wire NET_574;
wire NET_575;
wire NET_576;
wire NET_577;
wire NET_578;
wire NET_579;
wire NET_58;
wire NET_580;
wire NET_581;
wire NET_582;
wire NET_583;
wire NET_584;
wire NET_585;
wire NET_586;
wire NET_587;
wire NET_588;
wire NET_589;
wire NET_59;
wire NET_590;
wire NET_591;
wire NET_592;
wire NET_593;
wire NET_594;
wire NET_595;
wire NET_596;
wire NET_597;
wire NET_598;
wire NET_599;
wire NET_6;
wire NET_60;
wire NET_600;
wire NET_601;
wire NET_602;
wire NET_603;
wire NET_604;
wire NET_605;
wire NET_606;
wire NET_607;
wire NET_608;
wire NET_609;
wire NET_61;
wire NET_610;
wire NET_611;
wire NET_612;
wire NET_613;
wire NET_614;
wire NET_615;
wire NET_616;
wire NET_617;
wire NET_618;
wire NET_619;
wire NET_62;
wire NET_620;
wire NET_621;
wire NET_622;
wire NET_623;
wire NET_624;
wire NET_625;
wire NET_626;
wire NET_627;
wire NET_628;
wire NET_629;
wire NET_63;
wire NET_630;
wire NET_631;
wire NET_632;
wire NET_633;
wire NET_634;
wire NET_635;
wire NET_636;
wire NET_637;
wire NET_638;
wire NET_639;
wire NET_64;
wire NET_640;
wire NET_641;
wire NET_642;
wire NET_643;
wire NET_644;
wire NET_645;
wire NET_646;
wire NET_647;
wire NET_648;
wire NET_649;
wire NET_65;
wire NET_650;
wire NET_651;
wire NET_652;
wire NET_653;
wire NET_654;
wire NET_655;
wire NET_656;
wire NET_657;
wire NET_658;
wire NET_659;
wire NET_66;
wire NET_660;
wire NET_661;
wire NET_662;
wire NET_663;
wire NET_664;
wire NET_665;
wire NET_666;
wire NET_667;
wire NET_668;
wire NET_669;
wire NET_67;
wire NET_670;
wire NET_671;
wire NET_672;
wire NET_673;
wire NET_674;
wire NET_675;
wire NET_676;
wire NET_677;
wire NET_678;
wire NET_679;
wire NET_68;
wire NET_680;
wire NET_681;
wire NET_682;
wire NET_683;
wire NET_684;
wire NET_685;
wire NET_686;
wire NET_687;
wire NET_688;
wire NET_689;
wire NET_69;
wire NET_690;
wire NET_691;
wire NET_692;
wire NET_693;
wire NET_694;
wire NET_695;
wire NET_696;
wire NET_697;
wire NET_698;
wire NET_699;
wire NET_7;
wire NET_70;
wire NET_700;
wire NET_701;
wire NET_702;
wire NET_703;
wire NET_704;
wire NET_705;
wire NET_706;
wire NET_707;
wire NET_708;
wire NET_709;
wire NET_71;
wire NET_710;
wire NET_711;
wire NET_712;
wire NET_713;
wire NET_714;
wire NET_715;
wire NET_716;
wire NET_717;
wire NET_718;
wire NET_719;
wire NET_72;
wire NET_720;
wire NET_721;
wire NET_722;
wire NET_723;
wire NET_724;
wire NET_725;
wire NET_726;
wire NET_727;
wire NET_728;
wire NET_729;
wire NET_73;
wire NET_730;
wire NET_731;
wire NET_732;
wire NET_733;
wire NET_734;
wire NET_735;
wire NET_736;
wire NET_737;
wire NET_738;
wire NET_739;
wire NET_74;
wire NET_740;
wire NET_741;
wire NET_742;
wire NET_743;
wire NET_744;
wire NET_745;
wire NET_746;
wire NET_747;
wire NET_748;
wire NET_749;
wire NET_75;
wire NET_750;
wire NET_751;
wire NET_752;
wire NET_753;
wire NET_754;
wire NET_755;
wire NET_756;
wire NET_757;
wire NET_758;
wire NET_759;
wire NET_76;
wire NET_760;
wire NET_761;
wire NET_762;
wire NET_77;
wire NET_78;
wire NET_79;
wire NET_7_CAND3_TRSBL_17_tpGCLKBUF;
wire NET_7_CAND3_TRSBL_18_tpGCLKBUF;
wire NET_7_CAND3_TRSBL_19_tpGCLKBUF;
wire NET_7_CAND3_TRSBL_20_tpGCLKBUF;
wire NET_7_CAND3_TRSBL_21_tpGCLKBUF;
wire NET_7_CAND3_TRSBL_22_tpGCLKBUF;
wire NET_7_SQMUX_TRSBL3_tpGCLKBUF;
wire NET_8;
wire NET_80;
wire NET_81;
wire NET_82;
wire NET_83;
wire NET_83_CAND2_BRSTL_18_tpGCLKBUF;
wire NET_83_CAND2_BRSTL_19_tpGCLKBUF;
wire NET_83_CAND2_BRSTL_20_tpGCLKBUF;
wire NET_83_SQMUX_BRSTL2_tpGCLKBUF;
wire NET_84;
wire NET_85;
wire NET_86;
wire NET_87;
wire NET_88;
wire NET_89;
wire NET_9;
wire NET_90;
wire NET_91;
wire NET_92;
wire NET_93;
wire NET_94;
wire NET_95;
wire NET_96;
wire NET_97;
wire NET_98;
wire NET_99;
wire lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF;
wire lint_ADDR_int_13__CAND4_TLSTR_11_tpGCLKBUF;
wire lint_ADDR_int_13__CAND4_TLSTR_12_tpGCLKBUF;
wire lint_ADDR_int_13__CAND4_TLSTR_13_tpGCLKBUF;
wire lint_ADDR_int_13__CAND4_TLSTR_14_tpGCLKBUF;
wire lint_ADDR_int_13__CAND4_TLSTR_15_tpGCLKBUF;
wire lint_ADDR_int_13__SQMUX_TLSTR4_tpGCLKBUF;
wire lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF;
wire lint_ADDR_int_14__CAND5_TLSTR_11_tpGCLKBUF;
wire lint_ADDR_int_14__CAND5_TLSTR_12_tpGCLKBUF;
wire lint_ADDR_int_14__CAND5_TLSTR_13_tpGCLKBUF;
wire lint_ADDR_int_14__CAND5_TLSTR_14_tpGCLKBUF;
wire lint_ADDR_int_14__SQMUX_TLSTR5_tpGCLKBUF;
wire lint_GNT;
wire lint_GNT_dup_0;
wire lint_REQ;
wire lint_REQ_int;
wire lint_VALID;
wire lint_VALID_dup_0;
wire lint_WEN;
wire lint_WEN_int;
wire m0_coef_powerdn;
wire m0_coef_rclk;
wire m0_coef_wclk;
wire m0_coef_wdsel;
wire m0_coef_wdsel_dup_0;
wire m0_coef_we;
wire m0_coef_we_dup_0;
wire m0_m0_clk;
wire m0_m0_clken;
wire m0_m0_clken_dup_0;
wire m0_m0_clr;
wire m0_m0_clr_dup_0;
wire m0_m0_csel;
wire m0_m0_csel_dup_0;
wire m0_m0_osel;
wire m0_m0_osel_dup_0;
wire m0_m0_reset;
wire m0_m0_reset_dup_0;
wire m0_m0_rnd;
wire m0_m0_rnd_dup_0;
wire m0_m0_sat;
wire m0_m0_sat_dup_0;
wire m0_m0_tc;
wire m0_m0_tc_dup_0;
wire m0_m1_clk;
wire m0_m1_clken;
wire m0_m1_clken_dup_0;
wire m0_m1_clr;
wire m0_m1_clr_dup_0;
wire m0_m1_csel;
wire m0_m1_csel_dup_0;
wire m0_m1_osel;
wire m0_m1_osel_dup_0;
wire m0_m1_reset;
wire m0_m1_reset_dup_0;
wire m0_m1_rnd;
wire m0_m1_rnd_dup_0;
wire m0_m1_sat;
wire m0_m1_sat_dup_0;
wire m0_m1_tc;
wire m0_m1_tc_dup_0;
wire m0_oper0_powerdn;
wire m0_oper0_rclk;
wire m0_oper0_wclk;
wire m0_oper0_wdsel;
wire m0_oper0_wdsel_dup_0;
wire m0_oper0_we;
wire m0_oper0_we_dup_0;
wire m0_oper1_powerdn;
wire m0_oper1_rclk;
wire m0_oper1_wclk;
wire m0_oper1_wdsel;
wire m0_oper1_wdsel_dup_0;
wire m0_oper1_we;
wire m0_oper1_we_dup_0;
wire m1_coef_powerdn;
wire m1_coef_rclk;
wire m1_coef_wclk;
wire m1_coef_wdsel;
wire m1_coef_we;
wire m1_coef_we_dup_0;
wire m1_m0_clk;
wire m1_m0_clken;
wire m1_m0_clken_dup_0;
wire m1_m0_clr;
wire m1_m0_clr_dup_0;
wire m1_m0_csel;
wire m1_m0_csel_dup_0;
wire m1_m0_osel;
wire m1_m0_osel_dup_0;
wire m1_m0_reset;
wire m1_m0_reset_dup_0;
wire m1_m0_rnd;
wire m1_m0_rnd_dup_0;
wire m1_m0_sat;
wire m1_m0_sat_dup_0;
wire m1_m0_tc;
wire m1_m0_tc_dup_0;
wire m1_m1_clk;
wire m1_m1_clken;
wire m1_m1_clken_dup_0;
wire m1_m1_clr;
wire m1_m1_clr_dup_0;
wire m1_m1_csel;
wire m1_m1_csel_dup_0;
wire m1_m1_osel;
wire m1_m1_osel_dup_0;
wire m1_m1_reset;
wire m1_m1_reset_dup_0;
wire m1_m1_rnd;
wire m1_m1_rnd_dup_0;
wire m1_m1_sat;
wire m1_m1_sat_dup_0;
wire m1_m1_tc;
wire m1_m1_tc_dup_0;
wire m1_oper0_powerdn;
wire m1_oper0_rclk;
wire m1_oper0_wclk;
wire m1_oper0_wdsel;
wire m1_oper0_we;
wire m1_oper0_we_dup_0;
wire m1_oper1_powerdn;
wire m1_oper1_rclk;
wire m1_oper1_wclk;
wire m1_oper1_wdsel;
wire m1_oper1_we;
wire m1_oper1_we_dup_0;
wire not_RESET_0;
wire not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBL_17_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBL_18_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBL_23_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBL_24_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTL_17_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTL_18_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTL_22_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTR_28_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF;
wire not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTR_12_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF;
wire not_RESET_0_CAND3_TLSTR_9_tpGCLKBUF;
wire not_RESET_0_QMUX_BL1_tpGCLKBUF;
wire not_RESET_0_QMUX_BR1_tpGCLKBUF;
wire not_RESET_0_QMUX_TL3_tpGCLKBUF;
wire not_RESET_0_QMUX_TR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSBL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSBL3_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSBR3_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSTL3_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSTR3_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF;
wire not_RESET_1;
wire not_RESET_2;
wire not_RESET_3;
wire not_apb_fsm_0;
wire not_apb_fsm_1;
wire nx10146z1;
wire nx10146z2;
wire nx10775z1;
wire nx11310z2;
wire nx11311z2;
wire nx11312z2;
wire nx11313z3;
wire nx14650z1;
wire nx14650z1_CAND2_BRSBL_17_tpGCLKBUF;
wire nx14650z1_CAND2_BRSBL_18_tpGCLKBUF;
wire nx14650z1_SQMUX_BRSBL2_tpGCLKBUF;
wire nx15998z1;
wire nx15998z1_CAND2_TLSTR_13_tpGCLKBUF;
wire nx15998z1_CAND2_TLSTR_14_tpGCLKBUF;
wire nx15998z1_CAND2_TLSTR_15_tpGCLKBUF;
wire nx15998z1_CAND2_TLSTR_16_tpGCLKBUF;
wire nx15998z1_SQMUX_TLSTR2_tpGCLKBUF;
wire nx16907z1;
wire nx18281z1;
wire nx18281z1_CAND5_TRSTR_28_tpGCLKBUF;
wire nx18281z1_CAND5_TRSTR_29_tpGCLKBUF;
wire nx18281z1_SQMUX_TRSTR5_tpGCLKBUF;
wire nx19726z1;
wire nx19726z1_CAND2_BLSTR_10_tpGCLKBUF;
wire nx19726z1_CAND2_BLSTR_11_tpGCLKBUF;
wire nx19726z1_CAND2_BLSTR_12_tpGCLKBUF;
wire nx19726z1_CAND2_BLSTR_13_tpGCLKBUF;
wire nx19726z1_CAND2_BLSTR_14_tpGCLKBUF;
wire nx19726z1_CAND2_BLSTR_9_tpGCLKBUF;
wire nx19726z1_SQMUX_BLSTR2_tpGCLKBUF;
wire nx22245z1;
wire nx22245z1_CAND4_BLSBL_3_tpGCLKBUF;
wire nx22245z1_CAND4_BLSBL_4_tpGCLKBUF;
wire nx22245z1_CAND4_BLSBL_5_tpGCLKBUF;
wire nx22245z1_CAND4_BLSBL_6_tpGCLKBUF;
wire nx22245z1_CAND4_BLSBL_7_tpGCLKBUF;
wire nx22245z1_SQMUX_BLSBL4_tpGCLKBUF;
wire nx23147z1;
wire nx2520z1;
wire nx2520z1_CAND2_BRSBR_30_tpGCLKBUF;
wire nx2520z1_CAND2_BRSBR_31_tpGCLKBUF;
wire nx2520z1_CAND2_BRSBR_32_tpGCLKBUF;
wire nx2520z1_CAND2_BRSTR_30_tpGCLKBUF;
wire nx2520z1_CAND2_BRSTR_31_tpGCLKBUF;
wire nx2520z1_CAND2_BRSTR_32_tpGCLKBUF;
wire nx2520z1_QMUX_BR2_tpGCLKBUF;
wire nx2520z1_SQMUX_BRSBR2_tpGCLKBUF;
wire nx2520z1_SQMUX_BRSTR2_tpGCLKBUF;
wire nx25326z1;
wire nx25587z1;
wire nx25587z1_CAND2_TRSTR_25_tpGCLKBUF;
wire nx25587z1_CAND2_TRSTR_26_tpGCLKBUF;
wire nx25587z1_CAND2_TRSTR_27_tpGCLKBUF;
wire nx25587z1_SQMUX_TRSTR2_tpGCLKBUF;
wire nx25788z1;
wire nx25788z1_CAND3_BRSBR_29_tpGCLKBUF;
wire nx25788z1_CAND3_BRSBR_30_tpGCLKBUF;
wire nx25788z1_CAND3_BRSBR_31_tpGCLKBUF;
wire nx25788z1_CAND3_BRSBR_32_tpGCLKBUF;
wire nx25788z1_SQMUX_BRSBR3_tpGCLKBUF;
wire nx28356z1;
wire nx30664z1;
wire nx30664z1_CAND5_BRSBR_25_tpGCLKBUF;
wire nx30664z1_CAND5_BRSBR_26_tpGCLKBUF;
wire nx30664z1_CAND5_BRSBR_27_tpGCLKBUF;
wire nx30664z1_SQMUX_BRSBR5_tpGCLKBUF;
wire nx30923z1;
wire nx30923z1_CAND4_BRSTR_29_tpGCLKBUF;
wire nx30923z1_CAND4_BRSTR_30_tpGCLKBUF;
wire nx30923z1_CAND4_BRSTR_31_tpGCLKBUF;
wire nx30923z1_CAND4_BRSTR_32_tpGCLKBUF;
wire nx30923z1_SQMUX_BRSTR4_tpGCLKBUF;
wire nx32231z1;
wire nx32231z1_CAND2_TRSTL_17_tpGCLKBUF;
wire nx32231z1_CAND2_TRSTL_18_tpGCLKBUF;
wire nx32231z1_SQMUX_TRSTL2_tpGCLKBUF;
wire nx33579z1;
wire nx33579z1_CAND2_BLSBR_13_tpGCLKBUF;
wire nx33579z1_CAND2_BLSBR_14_tpGCLKBUF;
wire nx33579z1_CAND2_BLSBR_15_tpGCLKBUF;
wire nx33579z1_CAND2_BLSBR_16_tpGCLKBUF;
wire nx33579z1_SQMUX_BLSBR2_tpGCLKBUF;
wire nx34006z2;
wire nx34006z2_CAND2_TLSTL_4_tpGCLKBUF;
wire nx34006z2_CAND2_TLSTL_5_tpGCLKBUF;
wire nx34006z2_CAND2_TLSTL_6_tpGCLKBUF;
wire nx34006z2_CAND2_TLSTL_7_tpGCLKBUF;
wire nx34006z2_SQMUX_TLSTL2_tpGCLKBUF;
wire nx34850z1;
wire nx34850z1_CAND5_TLSTL_7_tpGCLKBUF;
wire nx34850z1_CAND5_TLSTL_8_tpGCLKBUF;
wire nx34850z1_SQMUX_TLSTL5_tpGCLKBUF;
wire nx36058z1;
wire nx36058z1_CAND2_TRSBR_29_tpGCLKBUF;
wire nx36058z1_CAND2_TRSBR_30_tpGCLKBUF;
wire nx36058z1_CAND2_TRSBR_31_tpGCLKBUF;
wire nx36058z1_CAND2_TRSBR_32_tpGCLKBUF;
wire nx36058z1_SQMUX_TRSBR2_tpGCLKBUF;
wire nx39840z1;
wire nx39840z1_CAND4_TLSTL_3_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_4_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_5_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_6_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_7_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_8_tpGCLKBUF;
wire nx39840z1_SQMUX_TLSTL4_tpGCLKBUF;
wire nx40728z1;
wire nx41193z1;
wire nx41193z1_CAND3_TRSTR_29_tpGCLKBUF;
wire nx41193z1_CAND3_TRSTR_30_tpGCLKBUF;
wire nx41193z1_CAND3_TRSTR_31_tpGCLKBUF;
wire nx41193z1_CAND3_TRSTR_32_tpGCLKBUF;
wire nx41193z1_SQMUX_TRSTR3_tpGCLKBUF;
wire nx44608z1;
wire nx44608z1_CAND1_TLSTL_1_tpGCLKBUF;
wire nx44608z1_CAND1_TLSTL_2_tpGCLKBUF;
wire nx44608z1_CAND1_TLSTL_3_tpGCLKBUF;
wire nx44608z1_CAND1_TLSTL_5_tpGCLKBUF;
wire nx44608z1_SQMUX_TLSTL1_tpGCLKBUF;
wire nx47611z1;
wire nx47611z1_CAND4_TRSTR_30_tpGCLKBUF;
wire nx47611z1_CAND4_TRSTR_31_tpGCLKBUF;
wire nx47611z1_CAND4_TRSTR_32_tpGCLKBUF;
wire nx47611z1_SQMUX_TRSTR4_tpGCLKBUF;
wire nx4939z1;
wire nx4939z1_CAND4_BLSTL_5_tpGCLKBUF;
wire nx4939z1_CAND4_BLSTL_6_tpGCLKBUF;
wire nx4939z1_CAND4_BLSTL_7_tpGCLKBUF;
wire nx4939z1_CAND4_BLSTL_8_tpGCLKBUF;
wire nx4939z1_SQMUX_BLSTL4_tpGCLKBUF;
wire nx49808z64;
wire nx49808z64_CAND2_TLSBR_10_tpGCLKBUF;
wire nx49808z64_CAND2_TLSBR_11_tpGCLKBUF;
wire nx49808z64_CAND2_TLSBR_12_tpGCLKBUF;
wire nx49808z64_CAND2_TLSBR_13_tpGCLKBUF;
wire nx49808z64_CAND2_TLSBR_14_tpGCLKBUF;
wire nx49808z64_CAND2_TLSBR_9_tpGCLKBUF;
wire nx49808z64_SQMUX_TLSBR2_tpGCLKBUF;
wire nx49871z1;
wire nx52746z1;
wire nx52746z1_CAND3_TRSBR_29_tpGCLKBUF;
wire nx52746z1_CAND3_TRSBR_30_tpGCLKBUF;
wire nx52746z1_CAND3_TRSBR_31_tpGCLKBUF;
wire nx52746z1_CAND3_TRSBR_32_tpGCLKBUF;
wire nx52746z1_SQMUX_TRSBR3_tpGCLKBUF;
wire nx53524z1;
wire nx53672z1;
wire nx53672z1_CAND4_BRSBR_28_tpGCLKBUF;
wire nx53672z1_CAND4_BRSBR_29_tpGCLKBUF;
wire nx53672z1_SQMUX_BRSBR4_tpGCLKBUF;
wire nx57881z1;
wire nx57881z1_CAND3_BRSTR_30_tpGCLKBUF;
wire nx57881z1_CAND3_BRSTR_31_tpGCLKBUF;
wire nx57881z1_CAND3_BRSTR_32_tpGCLKBUF;
wire nx57881z1_SQMUX_BRSTR3_tpGCLKBUF;
wire nx58292z1;
wire nx60509z1;
wire nx60831z1;
wire nx60831z1_CAND3_BLSBL_7_tpGCLKBUF;
wire nx60831z1_CAND3_BLSBL_8_tpGCLKBUF;
wire nx60831z1_SQMUX_BLSBL3_tpGCLKBUF;
wire nx65467z1;
wire nx7012z2;
wire nx7012z3;
wire nx8488z1;
wire nx9707z1;
wire nx9707z1_CAND2_BLSBL_1_tpGCLKBUF;
wire nx9707z1_CAND2_BLSBL_2_tpGCLKBUF;
wire nx9707z1_CAND2_BLSBL_3_tpGCLKBUF;
wire nx9707z1_CAND2_BLSBL_5_tpGCLKBUF;
wire nx9707z1_CAND2_BLSTL_1_tpGCLKBUF;
wire nx9707z1_CAND2_BLSTL_3_tpGCLKBUF;
wire nx9707z1_CAND2_BLSTL_5_tpGCLKBUF;
wire nx9707z1_QMUX_BL2_tpGCLKBUF;
wire nx9707z1_SQMUX_BLSBL2_tpGCLKBUF;
wire nx9707z1_SQMUX_BLSTL2_tpGCLKBUF;
wire saved_REQ;
wire tcdm_clk_p0;
wire tcdm_clk_p1;
wire tcdm_clk_p2;
wire tcdm_clk_p3;
wire tcdm_gnt_p0;
wire tcdm_gnt_p0_int;
wire tcdm_gnt_p1;
wire tcdm_gnt_p1_int;
wire tcdm_gnt_p2;
wire tcdm_gnt_p2_int;
wire tcdm_gnt_p3;
wire tcdm_gnt_p3_int;
wire tcdm_req_p0;
wire tcdm_req_p0_dup_0;
wire tcdm_req_p1;
wire tcdm_req_p1_dup_0;
wire tcdm_req_p2;
wire tcdm_req_p2_dup_0;
wire tcdm_req_p3;
wire tcdm_req_p3_dup_0;
wire tcdm_valid_p0;
wire tcdm_valid_p0_int;
wire tcdm_valid_p0_int_CAND1_TLSBR_12_tpGCLKBUF;
wire tcdm_valid_p0_int_CAND1_TLSBR_13_tpGCLKBUF;
wire tcdm_valid_p0_int_CAND1_TLSBR_14_tpGCLKBUF;
wire tcdm_valid_p0_int_CAND1_TLSBR_15_tpGCLKBUF;
wire tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF;
wire tcdm_valid_p0_int_SQMUX_TLSBR1_tpGCLKBUF;
wire tcdm_valid_p1;
wire tcdm_valid_p1_int;
wire tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF;
wire tcdm_valid_p1_int_CAND5_TRSBL_18_tpGCLKBUF;
wire tcdm_valid_p1_int_CAND5_TRSBL_19_tpGCLKBUF;
wire tcdm_valid_p1_int_CAND5_TRSBL_20_tpGCLKBUF;
wire tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF;
wire tcdm_valid_p1_int_CAND5_TRSBL_22_tpGCLKBUF;
wire tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF;
wire tcdm_valid_p2;
wire tcdm_valid_p2_int;
wire tcdm_valid_p3;
wire tcdm_valid_p3_int;
wire tcdm_we_p0;
wire tcdm_we_p0_dup_0;
wire tcdm_we_p1;
wire tcdm_we_p1_dup_0;
wire tcdm_we_p2;
wire tcdm_we_p2_dup_0;
wire tcdm_we_p3;
wire tcdm_we_p3_dup_0;
wire [5:0] CLK;
wire [5:0] CLK_int;
wire [3:0] RESET;
wire [3:0] RESET_int;
wire [1:0] apb_fsm;
wire [2:0] cnt1;
wire [2:0] cnt2;
wire [2:0] cnt3;
wire [2:0] cnt4;
wire [2:0] cnt5;
wire [15:0] events_o;
wire [79:0] fpgaio_in;
wire [79:0] fpgaio_in_int;
wire [79:0] fpgaio_oe;
wire [79:0] fpgaio_oe_dup_0;
wire [79:0] fpgaio_out;
wire [79:0] fpgaio_out_dup_0;
wire [15:0] i_events;
wire [19:0] lint_ADDR;
wire [19:0] lint_ADDR_int;
wire [3:0] lint_BE;
wire [3:0] lint_BE_int;
wire [31:0] lint_RDATA;
wire [31:0] lint_RDATA_dup_0;
wire [31:0] lint_WDATA;
wire [31:0] lint_WDATA_int;
wire [11:0] m0_coef_raddr;
wire [11:0] m0_coef_raddr_dup_0;
wire [31:0] m0_coef_rdata;
wire [31:0] m0_coef_rdata_int;
wire [1:0] m0_coef_rmode;
wire [1:0] m0_coef_rmode_dup_0;
wire [11:0] m0_coef_waddr;
wire [11:0] m0_coef_waddr_dup_0;
wire [31:0] m0_coef_wdata;
wire [31:0] m0_coef_wdata_dup_0;
wire [1:0] m0_coef_wmode;
wire [1:0] m0_coef_wmode_dup_0;
wire [31:0] m0_m0_coef_in;
wire [30:7] m0_m0_control;
wire [31:0] m0_m0_dataout;
wire [31:0] m0_m0_dataout_int;
wire [1:0] m0_m0_mode;
wire [1:0] m0_m0_mode_dup_0;
wire [31:0] m0_m0_oper_in;
wire [5:0] m0_m0_outsel;
wire [5:0] m0_m0_outsel_dup_0;
wire [31:0] m0_m1_coef_in;
wire [30:7] m0_m1_control;
wire [31:0] m0_m1_dataout;
wire [31:0] m0_m1_dataout_int;
wire [1:0] m0_m1_mode;
wire [1:0] m0_m1_mode_dup_0;
wire [31:0] m0_m1_oper_in;
wire [5:0] m0_m1_outsel;
wire [5:0] m0_m1_outsel_dup_0;
wire [11:0] m0_oper0_raddr;
wire [11:0] m0_oper0_raddr_dup_0;
wire [31:0] m0_oper0_rdata;
wire [31:0] m0_oper0_rdata_int;
wire [1:0] m0_oper0_rmode;
wire [1:0] m0_oper0_rmode_dup_0;
wire [11:0] m0_oper0_waddr;
wire [11:0] m0_oper0_waddr_dup_0;
wire [31:0] m0_oper0_wdata;
wire [31:0] m0_oper0_wdata_dup_0;
wire [1:0] m0_oper0_wmode;
wire [1:0] m0_oper0_wmode_dup_0;
wire [11:0] m0_oper1_raddr;
wire [11:0] m0_oper1_raddr_dup_0;
wire [31:0] m0_oper1_rdata;
wire [31:0] m0_oper1_rdata_int;
wire [1:0] m0_oper1_rmode;
wire [1:0] m0_oper1_rmode_dup_0;
wire [11:0] m0_oper1_waddr;
wire [11:0] m0_oper1_waddr_dup_0;
wire [31:0] m0_oper1_wdata;
wire [31:0] m0_oper1_wdata_dup_0;
wire [1:0] m0_oper1_wmode;
wire [1:0] m0_oper1_wmode_dup_0;
wire [31:15] m0_ram_control;
wire [11:0] m1_coef_raddr;
wire [11:0] m1_coef_raddr_dup_0;
wire [31:0] m1_coef_rdata;
wire [31:0] m1_coef_rdata_int;
wire [1:0] m1_coef_rmode;
wire [11:0] m1_coef_waddr;
wire [11:0] m1_coef_waddr_dup_0;
wire [31:0] m1_coef_wdata;
wire [31:0] m1_coef_wdata_dup_0;
wire [1:0] m1_coef_wmode;
wire [31:0] m1_m0_coef_in;
wire [30:7] m1_m0_control;
wire [31:0] m1_m0_dataout;
wire [31:0] m1_m0_dataout_int;
wire [1:0] m1_m0_mode;
wire [1:0] m1_m0_mode_dup_0;
wire [31:0] m1_m0_oper_in;
wire [5:0] m1_m0_outsel;
wire [5:0] m1_m0_outsel_dup_0;
wire [31:0] m1_m1_coef_in;
wire [30:0] m1_m1_control;
wire [31:0] m1_m1_dataout;
wire [31:0] m1_m1_dataout_int;
wire [1:0] m1_m1_mode;
wire [1:0] m1_m1_mode_dup_0;
wire [31:0] m1_m1_oper_in;
wire [5:0] m1_m1_outsel;
wire [11:0] m1_oper0_raddr;
wire [11:0] m1_oper0_raddr_dup_0;
wire [31:0] m1_oper0_rdata;
wire [31:0] m1_oper0_rdata_int;
wire [1:0] m1_oper0_rmode;
wire [11:0] m1_oper0_waddr;
wire [11:0] m1_oper0_waddr_dup_0;
wire [31:0] m1_oper0_wdata;
wire [31:0] m1_oper0_wdata_dup_0;
wire [1:0] m1_oper0_wmode;
wire [11:0] m1_oper1_raddr;
wire [11:0] m1_oper1_raddr_dup_0;
wire [31:0] m1_oper1_rdata;
wire [31:0] m1_oper1_rdata_int;
wire [1:0] m1_oper1_rmode;
wire [11:0] m1_oper1_waddr;
wire [11:0] m1_oper1_waddr_dup_0;
wire [31:0] m1_oper1_wdata;
wire [31:0] m1_oper1_wdata_dup_0;
wire [1:0] m1_oper1_wmode;
wire [31:0] m1_ram_control;
wire [19:0] tcdm_addr_p0;
wire [19:0] tcdm_addr_p0_dup_0;
wire [19:0] tcdm_addr_p1;
wire [19:0] tcdm_addr_p1_dup_0;
wire [19:0] tcdm_addr_p2;
wire [19:0] tcdm_addr_p2_dup_0;
wire [19:0] tcdm_addr_p3;
wire [19:0] tcdm_addr_p3_dup_0;
wire [3:0] tcdm_be_p0;
wire [3:0] tcdm_be_p0_dup_0;
wire [3:0] tcdm_be_p1;
wire [3:0] tcdm_be_p1_dup_0;
wire [3:0] tcdm_be_p2;
wire [3:0] tcdm_be_p2_dup_0;
wire [3:0] tcdm_be_p3;
wire [3:0] tcdm_be_p3_dup_0;
wire [31:0] tcdm_rdata_p0;
wire [31:0] tcdm_rdata_p0_int;
wire [31:0] tcdm_rdata_p1;
wire [31:0] tcdm_rdata_p1_int;
wire [31:0] tcdm_rdata_p2;
wire [31:0] tcdm_rdata_p2_int;
wire [31:0] tcdm_rdata_p3;
wire [31:0] tcdm_rdata_p3_int;
wire [31:0] tcdm_result_p0;
wire [31:0] tcdm_result_p1;
wire [31:0] tcdm_result_p2;
wire [31:0] tcdm_result_p3;
wire [31:0] tcdm_wdata_p0;
wire [31:0] tcdm_wdata_p0_dup_0;
wire [31:0] tcdm_wdata_p1;
wire [31:0] tcdm_wdata_p1_dup_0;
wire [31:0] tcdm_wdata_p2;
wire [31:0] tcdm_wdata_p2_dup_0;
wire [31:0] tcdm_wdata_p3;
wire [31:0] tcdm_wdata_p3_dup_0;

	LOGIC_0 QL_INST_A3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[13]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A8_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_in_int[31]),.B0I1(fpgaio_oe_dup_0[31]),.B0I2(NET_64),.B0I3(NET_30),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_in_int[31]),.T0I1(fpgaio_oe_dup_0[31]),.T0I2(NET_64),.T0I3(NET_30),.TB0S(NET_8),.C0Z(NET_613),.Q0Z(fpgaio_oe_dup_0[31]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A8_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(fpgaio_in_int[20]),.B1I1(NET_30),.B1I2(NET_64),.B1I3(fpgaio_oe_dup_0[20]),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.T1I0(NET_64),.T1I1(fpgaio_oe_dup_0[20]),.T1I2(fpgaio_in_int[20]),.T1I3(NET_30),.TB1S(NET_8),.C1Z(NET_397),.Q1Z(fpgaio_oe_dup_0[30]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_A8_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B2I0(fpgaio_oe_dup_0[16]),.B2I1(fpgaio_in_int[16]),.B2I2(NET_64),.B2I3(NET_30),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_oe_dup_0[16]),.T2I1(fpgaio_in_int[16]),.T2I2(NET_64),.T2I3(NET_30),.TB2S(NET_8),.C2Z(NET_323),.Q2Z(fpgaio_oe_dup_0[27]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_A8_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B3I0(NET_64),.B3I1(NET_30),.B3I2(fpgaio_in_int[25]),.B3I3(fpgaio_oe_dup_0[25]),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_in_int[25]),.T3I1(fpgaio_oe_dup_0[25]),.T3I2(NET_64),.T3I3(NET_30),.TB3S(NET_8),.C3Z(NET_507),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_A9_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_in_int[30]),.B0I1(NET_30),.B0I2(NET_64),.B0I3(fpgaio_oe_dup_0[30]),.T0I0(fpgaio_in_int[30]),.T0I1(NET_30),.T0I2(NET_64),.T0I3(fpgaio_oe_dup_0[30]),.TB0S(NET_8),.C0Z(NET_595),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_A9_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B1I0(NET_10),.B1I1(fpgaio_in_int[5]),.B1I2(NET_8),.B1I3(fpgaio_in_int[37]),.T1I0(NET_8),.T1I1(fpgaio_in_int[37]),.T1I2(NET_10),.T1I3(fpgaio_in_int[5]),.TB1S(NET_64),.C1Z(NET_661),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_A9_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_8),.B2I1(fpgaio_in_int[35]),.B2I2(NET_10),.B2I3(fpgaio_in_int[3]),.T2I0(NET_8),.T2I1(fpgaio_in_int[35]),.T2I2(NET_10),.T2I3(fpgaio_in_int[3]),.TB2S(NET_64),.C2Z(NET_700),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_A9_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B3I0(fpgaio_oe_dup_0[27]),.B3I1(NET_64),.B3I2(NET_30),.B3I3(fpgaio_in_int[27]),.T3I0(NET_30),.T3I1(fpgaio_in_int[27]),.T3I2(fpgaio_oe_dup_0[27]),.T3I3(NET_64),.TB3S(NET_8),.C3Z(NET_542),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_A10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A10_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B2I0(fpgaio_in_int[15]),.B2I1(NET_10),.B2I2(NET_8),.B2I3(fpgaio_in_int[47]),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[15]),.T2I1(NET_10),.T2I2(NET_8),.T2I3(fpgaio_in_int[47]),.TB2S(NET_64),.C2Z(NET_306),.Q2Z(fpgaio_oe_dup_0[29]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_A10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A13_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B1I0(fpgaio_in_int[42]),.B1I1(NET_10),.B1I2(NET_8),.B1I3(fpgaio_in_int[10]),.T1I0(NET_8),.T1I1(fpgaio_in_int[10]),.T1I2(fpgaio_in_int[42]),.T1I3(NET_10),.TB1S(NET_64),.C1Z(NET_188),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_A13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A13_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B3I0(NET_10),.B3I1(fpgaio_in_int[45]),.B3I2(NET_8),.B3I3(fpgaio_in_int[13]),.T3I0(NET_8),.T3I1(fpgaio_in_int[13]),.T3I2(NET_10),.T3I3(fpgaio_in_int[45]),.TB3S(NET_64),.C3Z(NET_247),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_A14_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_8),.B0I1(fpgaio_in_int[40]),.B0I2(fpgaio_in_int[8]),.B0I3(NET_10),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(NET_8),.T0I1(fpgaio_in_int[40]),.T0I2(fpgaio_in_int[8]),.T0I3(NET_10),.TB0S(NET_64),.C0Z(NET_287),.Q0Z(fpgaio_oe_dup_0[21]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A14_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B3I0(fpgaio_in_int[9]),.B3I1(NET_10),.B3I2(NET_8),.B3I3(fpgaio_in_int[41]),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.T3I0(NET_8),.T3I1(fpgaio_in_int[41]),.T3I2(fpgaio_in_int[9]),.T3I3(NET_10),.TB3S(NET_64),.C3Z(NET_166),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_A15_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_in_int[14]),.B0I1(fpgaio_in_int[46]),.B0I2(NET_8),.B0I3(NET_10),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_in_int[14]),.T0I1(fpgaio_in_int[46]),.T0I2(NET_8),.T0I3(NET_10),.TB0S(NET_64),.C0Z(NET_267),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A15_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(fpgaio_in_int[43]),.B1I1(fpgaio_in_int[11]),.B1I2(NET_10),.B1I3(NET_8),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.T1I0(NET_10),.T1I1(NET_8),.T1I2(fpgaio_in_int[43]),.T1I3(fpgaio_in_int[11]),.TB1S(NET_64),.C1Z(NET_207),.Q1Z(fpgaio_oe_dup_0[17]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_A15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A16_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(fpgaio_oe_dup_0[18]),.T1I1(NET_123),.T1I2(fpgaio_oe_dup_0[50]),.T1I3(NET_126),.TB1S(GND),.C1Z(NET_358),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_A16_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.T2I0(fpgaio_oe_dup_0[17]),.T2I1(NET_123),.T2I2(fpgaio_oe_dup_0[49]),.T2I3(NET_126),.TB2S(GND),.C2Z(NET_340),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_A16_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(fpgaio_oe_dup_0[51]),.T3I1(NET_123),.T3I2(fpgaio_oe_dup_0[19]),.T3I3(NET_126),.TB3S(GND),.C3Z(NET_377),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_A17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_126),.B0I1(fpgaio_oe_dup_0[28]),.B0I2(fpgaio_oe_dup_0[60]),.B0I3(NET_123),.B0Z(NET_558),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A17_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_126),.T1I1(fpgaio_oe_dup_0[29]),.T1I2(fpgaio_oe_dup_0[61]),.T1I3(NET_123),.TB1S(GND),.C1Z(NET_576),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_A17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A18_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001000000000000),.B0I0(lint_ADDR_int[11]),.B0I1(GND),.B0I2(NET_10),.B0I3(NET_30),.T0I0(fpgaio_oe_dup_0[24]),.T0I1(NET_126),.T0I2(NET_123),.T0I3(fpgaio_oe_dup_0[56]),.TB0S(GND),.B0Z(NET_126),.C0Z(NET_488),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_A18_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(fpgaio_oe_dup_0[23]),.T1I1(fpgaio_oe_dup_0[55]),.T1I2(NET_123),.T1I3(NET_126),.TB1S(GND),.C1Z(NET_449),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_A18_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B2I0(fpgaio_oe_dup_0[54]),.B2I1(NET_126),.B2I2(NET_123),.B2I3(fpgaio_oe_dup_0[22]),.T2I0(fpgaio_oe_dup_0[26]),.T2I1(fpgaio_oe_dup_0[58]),.T2I2(NET_123),.T2I3(NET_126),.TB2S(GND),.B2Z(NET_431),.C2Z(NET_523),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_A18_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(fpgaio_oe_dup_0[53]),.T3I1(fpgaio_oe_dup_0[21]),.T3I2(NET_123),.T3I3(NET_126),.TB3S(GND),.C3Z(NET_413),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_A19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[56]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[53]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[51]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(fpgaio_in_int[57]),.B1I1(NET_322),.B1I2(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.B1I3(fpgaio_oe_dup_0[57]),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T1I0(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.T1I1(fpgaio_oe_dup_0[57]),.T1I2(fpgaio_in_int[57]),.T1I3(NET_322),.TB1S(NET_507),.C1Z(NET_505),.Q1Z(fpgaio_oe_dup_0[49]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_A20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(fpgaio_in_int[59]),.B2I1(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.B2I2(fpgaio_oe_dup_0[59]),.B2I3(NET_322),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[59]),.T2I1(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.T2I2(fpgaio_oe_dup_0[59]),.T2I3(NET_322),.TB2S(NET_542),.C2Z(NET_540),.Q2Z(fpgaio_oe_dup_0[59]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_A20_3 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_10),.T3I2(GND),.T3I3(NET_64),.TB3S(GND),.C3Z(NET_322),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_A21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.B0I1(NET_322),.B0I2(fpgaio_oe_dup_0[63]),.B0I3(fpgaio_in_int[63]),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T0I0(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.T0I1(NET_322),.T0I2(fpgaio_oe_dup_0[63]),.T0I3(fpgaio_in_int[63]),.TB0S(NET_613),.C0Z(NET_611),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[23]),.Q2EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[55]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[58]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_322),.B0I1(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.B0I2(fpgaio_in_int[48]),.B0I3(fpgaio_oe_dup_0[48]),.CD0S(VCC),.Q0DI(lint_WDATA_int[28]),.Q0EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T0I0(NET_322),.T0I1(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.T0I2(fpgaio_in_int[48]),.T0I3(fpgaio_oe_dup_0[48]),.TB0S(NET_323),.C0Z(NET_320),.Q0Z(fpgaio_oe_dup_0[60]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[63]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_322),.B2I1(fpgaio_in_int[52]),.B2I2(fpgaio_oe_dup_0[52]),.B2I3(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(NET_322),.T2I1(fpgaio_in_int[52]),.T2I2(fpgaio_oe_dup_0[52]),.T2I3(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.TB2S(NET_397),.C2Z(NET_395),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_A22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(fpgaio_in_int[62]),.B3I1(fpgaio_oe_dup_0[62]),.B3I2(NET_322),.B3I3(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T3I0(NET_322),.T3I1(NET_29_CAND5_BLSTL_1_tpGCLKBUF),.T3I2(fpgaio_in_int[62]),.T3I3(fpgaio_oe_dup_0[62]),.TB3S(NET_595),.C3Z(NET_593),.Q3Z(fpgaio_oe_dup_0[40]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_A23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[52]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[45]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[54]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[57]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[62]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[61]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[50]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A25_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_127),.B0I1(fpgaio_in_int[32]),.B0I2(fpgaio_oe_dup_0[32]),.B0I3(NET_126),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(NET_127),.T0I1(fpgaio_in_int[34]),.T0I2(fpgaio_oe_dup_0[34]),.T0I3(NET_126),.TB0S(GND),.B0Z(NET_122),.C0Z(NET_724),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[48]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[32]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[34]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A26_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(NET_126),.T0I1(fpgaio_oe_dup_0[38]),.T0I2(NET_127),.T0I3(fpgaio_in_int[38]),.TB0S(GND),.C0Z(NET_643),.Q0Z(fpgaio_oe_dup_0[38]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[39]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_126),.B2I1(fpgaio_oe_dup_0[44]),.B2I2(NET_127),.B2I3(fpgaio_in_int[44]),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.B2Z(NET_231),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A26_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.T3I0(NET_126),.T3I1(fpgaio_in_int[39]),.T3I2(NET_127),.T3I3(fpgaio_oe_dup_0[39]),.C3Z(NET_477),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_B3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx44608z1_CAND1_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx44608z1_CAND1_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx44608z1_CAND1_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx44608z1_CAND1_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B9_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_in_int[36]),.B0I1(NET_8),.B0I2(NET_10),.B0I3(fpgaio_in_int[4]),.T0I0(fpgaio_in_int[36]),.T0I1(NET_8),.T0I2(NET_10),.T0I3(fpgaio_in_int[4]),.TB0S(NET_64),.C0Z(NET_681),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_B9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B9_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B3I0(NET_10),.B3I1(fpgaio_in_int[1]),.B3I2(fpgaio_in_int[33]),.B3I3(NET_8),.T3I0(fpgaio_in_int[33]),.T3I1(NET_8),.T3I2(NET_10),.T3I3(fpgaio_in_int[1]),.TB3S(NET_64),.C3Z(NET_53),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_B18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B2I0(NET_8),.B2I1(lint_ADDR_int[11]),.B2I2(GND),.B2I3(NET_30),.B2Z(NET_123),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B0I0(NET_10),.B0I1(GND),.B0I2(GND),.B0I3(NET_30),.B0Z(NET_29),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx9707z1_CAND2_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[44]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx9707z1_CAND2_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[47]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx9707z1_CAND2_BLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[46]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx44608z1_CAND1_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx44608z1_CAND1_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx44608z1_CAND1_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx44608z1_CAND1_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx39840z1_CAND4_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx39840z1_CAND4_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx44608z1_CAND1_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[67]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[78]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C14_0 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.T0I0(NET_8),.T0I1(lint_ADDR_int[11]),.T0I2(GND),.T0I3(NET_64),.TB0S(GND),.C0Z(NET_111),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_C14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[71]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C17_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[5]),.T1I1(lint_ADDR_int[3]),.T1I2(lint_ADDR_int[6]),.T1I3(lint_ADDR_int[4]),.C1Z(NET_64),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_C17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C20_3 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_10),.T3I1(GND),.T3I2(NET_64),.T3I3(lint_ADDR_int[11]),.C3Z(NET_127),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_C21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx9707z1_CAND2_BLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[42]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx9707z1_CAND2_BLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[37]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx9707z1_CAND2_BLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[36]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx9707z1_CAND2_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[43]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx22245z1_CAND4_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[21]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx22245z1_CAND4_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx22245z1_CAND4_BLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_3_padClk),.QRT(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[25]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[29]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[27]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[20]),.Q2EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[20]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[69]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[8]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[72]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[68]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[79]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[77]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[64]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_129),.B0I1(NET_111),.B0I2(m1_m1_control[21]),.B0I3(fpgaio_in_int[21]),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.B0Z(NET_416),.Q0Z(m1_m1_control[26]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D15_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[21]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.T1I0(NET_129),.T1I1(NET_111),.T1I2(fpgaio_in_int[24]),.T1I3(m1_m1_control[24]),.C1Z(NET_491),.Q1Z(m1_m1_control[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_D15_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[26]),.T2I1(NET_111),.T2I2(NET_129),.T2I3(m1_m1_control[26]),.TB2S(GND),.C2Z(NET_526),.Q2Z(m1_m1_control[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_D15_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[24]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF),.QST(GND),.T3I0(NET_129),.T3I1(m1_m1_control[22]),.T3I2(fpgaio_in_int[22]),.T3I3(NET_111),.C3Z(NET_434),.Q3Z(m1_m1_control[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_D19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_GNT_dup_0),.Q0EN(not_apb_fsm_1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(lint_VALID_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D19_1 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[5]),.T1I1(lint_ADDR_int[4]),.T1I2(lint_ADDR_int[3]),.T1I3(lint_ADDR_int[6]),.C1Z(NET_30),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_D19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[24]),.Q3EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[22]),.Q0EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[20]),.Q3EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_4_padClk),.QRT(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[6]),.Q3EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_waddr_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[3]),.Q0EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_waddr_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx44608z1_CAND1_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx44608z1_CAND1_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx39840z1_CAND4_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx39840z1_CAND4_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx39840z1_CAND4_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E8_1 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(NET_30),.T1I2(NET_8),.T1I3(GND),.TB1S(GND),.C1Z(NET_58),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_E8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx44608z1_CAND1_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E9_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.T0I0(NET_123),.T0I1(fpgaio_oe_dup_0[7]),.T0I2(tcdm_rdata_p0_int[7]),.T0I3(NET_124),.TB0S(GND),.C0Z(NET_476),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E9_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[21]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.T1I0(NET_123),.T1I1(fpgaio_oe_dup_0[12]),.T1I2(NET_124),.T1I3(tcdm_rdata_p0_int[12]),.TB1S(GND),.C1Z(NET_230),.Q1Z(fpgaio_out_dup_0[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_E9_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_123),.B2I1(fpgaio_oe_dup_0[2]),.B2I2(tcdm_rdata_p0_int[2]),.B2I3(NET_124),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.T2I0(NET_123),.T2I1(fpgaio_oe_dup_0[0]),.T2I2(tcdm_rdata_p0_int[0]),.T2I3(NET_124),.TB2S(GND),.B2Z(NET_723),.C2Z(NET_121),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_E9_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.T3I0(NET_123),.T3I1(tcdm_rdata_p0_int[6]),.T3I2(NET_124),.T3I3(fpgaio_oe_dup_0[6]),.C3Z(NET_642),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_E10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[69]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[70]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[75]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[73]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[77]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[74]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[64]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[71]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[66]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[76]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[76]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_129),.B0I1(NET_111),.B0I2(fpgaio_in_int[29]),.B0I3(m1_m1_control[29]),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.B0Z(NET_579),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E15_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.T1I0(NET_129),.T1I1(fpgaio_in_int[19]),.T1I2(m1_m1_control[19]),.T1I3(NET_111),.C1Z(NET_380),.Q1Z(m1_m1_control[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_E15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_129),.B2I1(fpgaio_in_int[23]),.B2I2(m1_m1_control[23]),.B2I3(NET_111),.CD2S(VCC),.Q2DI(lint_WDATA_int[23]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.B2Z(NET_452),.Q2Z(m1_m1_control[23]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_control[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E16_0 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0000100000000000),.B0I0(NET_122),.B0I1(NET_120),.B0I2(GND),.B0I3(NET_121),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(NET_642),.T0I2(NET_641),.T0I3(NET_643),.TB0S(GND),.B0Z(NET_78),.C0Z(NET_624),.Q0Z(m1_m1_control[0]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(NET_129),.B1I1(m1_m1_control[7]),.B1I2(fpgaio_out_dup_0[71]),.B1I3(NET_128),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[71]),.T1I1(NET_128),.T1I2(NET_129),.T1I3(m1_m1_control[7]),.TB1S(NET_478),.C1Z(NET_475),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_E16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_m1_control[0]),.B2I1(NET_128),.B2I2(NET_129),.B2I3(fpgaio_out_dup_0[64]),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.T2I0(m1_m1_control[0]),.T2I1(NET_128),.T2I2(NET_129),.T2I3(fpgaio_out_dup_0[64]),.TB2S(NET_130),.C2Z(NET_120),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_E16_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF),.QST(GND),.T3I0(NET_477),.T3I1(GND),.T3I2(NET_476),.T3I3(NET_475),.C3Z(NET_458),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_E17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(fpgaio_out_dup_0[66]),.B1I1(NET_128),.B1I2(m1_m1_control[2]),.B1I3(NET_129),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_control[2]),.T1I1(NET_129),.T1I2(fpgaio_out_dup_0[66]),.T1I3(NET_128),.TB1S(NET_725),.C1Z(NET_722),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_E17_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T2I0(NET_724),.T2I1(NET_723),.T2I2(NET_722),.T2I3(GND),.TB2S(GND),.C2Z(NET_705),.Q2Z(m1_m1_control[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_E17_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(NET_229),.T3I1(NET_230),.T3I2(NET_231),.T3I3(GND),.C3Z(NET_212),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_E18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_488),.B0I1(NET_490),.B0I2(NET_491),.B0I3(NET_489),.T0I0(NET_488),.T0I1(NET_490),.T0I2(NET_491),.T0I3(NET_489),.TB0S(NET_492),.C0Z(NET_480),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_E18_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(GND),.T1I1(RESET_int[3]),.T1I2(GND),.T1I3(GND),.TB1S(GND),.C1Z(not_RESET_3),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_E18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_416),.B2I1(NET_414),.B2I2(NET_415),.B2I3(NET_413),.T2I0(NET_416),.T2I1(NET_414),.T2I2(NET_415),.T2I3(NET_413),.TB2S(NET_417),.C2Z(NET_405),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_E18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_450),.B3I1(NET_452),.B3I2(NET_449),.B3I3(NET_451),.T3I0(NET_449),.T3I1(NET_451),.T3I2(NET_450),.T3I3(NET_452),.TB3S(NET_453),.C3Z(NET_441),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_E19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E19_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx4939z1_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(NET_602),.T1I1(GND),.T1I2(NET_67),.T1I3(GND),.TB1S(GND),.C1Z(nx9707z1),.Q1Z(fpgaio_out_dup_0[35]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_E19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx4939z1_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[41]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E20_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_in_int[54]),.T1I1(NET_127),.T1I2(m1_m0_control[22]),.T1I3(NET_119),.TB1S(GND),.C1Z(NET_435),.Q1Z(m1_m0_control[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_E20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx4939z1_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[53]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E20_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_in_int[55]),.T3I1(NET_127),.T3I2(m1_m0_control[23]),.T3I3(NET_119),.C3Z(NET_453),.Q3Z(m1_m0_control[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_E21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(fpgaio_in_int[53]),.B0I1(NET_127),.B0I2(m1_m0_control[21]),.B0I3(NET_119),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0Z(NET_417),.Q0Z(m1_m0_control[19]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx4939z1_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[44]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_119),.B2I1(NET_127),.B2I2(m1_m0_control[24]),.B2I3(fpgaio_in_int[56]),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B2Z(NET_492),.Q2Z(m1_m0_control[21]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E21_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[24]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(NET_119),.T3I1(NET_127),.T3I2(fpgaio_in_int[51]),.T3I3(m1_m0_control[19]),.C3Z(NET_381),.Q3Z(m1_m0_control[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_E22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx4939z1_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[32]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx4939z1_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[36]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx9707z1_CAND2_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[35]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E23_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_in_int[61]),.T0I1(m1_m0_control[29]),.T0I2(NET_119),.T0I3(NET_127),.TB0S(GND),.C0Z(NET_580),.Q0Z(m1_m0_control[29]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx4939z1_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[62]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx4939z1_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[57]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx4939z1_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[52]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx9707z1_CAND2_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[33]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[9]),.Q1EN(nx9707z1_CAND2_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[41]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[2]),.Q3EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_waddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[8]),.Q0EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_waddr_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[9]),.Q1EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_waddr_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[5]),.Q0EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_waddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[4]),.Q1EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_waddr_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[1]),.Q2EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_waddr_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[9]),.Q3EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_waddr_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[8]),.Q0EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_waddr_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[2]),.Q1EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_waddr_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[7]),.Q3EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_waddr_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_wdata_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_wdata_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_waddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_wdata_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdata_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx39840z1_CAND4_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[68]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[74]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[65]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[75]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_20),.B0I1(fpgaio_oe_dup_0[74]),.B0I2(i_events[10]),.B0I3(NET_21),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.B0Z(NET_174),.Q0Z(i_events[8]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(i_events[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F12_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_20),.B2I1(NET_21),.B2I2(fpgaio_oe_dup_0[73]),.B2I3(i_events[9]),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.T2I0(NET_20),.T2I1(fpgaio_oe_dup_0[69]),.T2I2(i_events[5]),.T2I3(NET_21),.TB2S(GND),.B2Z(NET_152),.C2Z(NET_647),.Q2Z(i_events[5]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_F12_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(NET_20),.T3I1(i_events[8]),.T3I2(fpgaio_oe_dup_0[72]),.T3I3(NET_21),.TB3S(GND),.C3Z(NET_273),.Q3Z(i_events[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_F13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q0Z(i_events[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[70]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(fpgaio_oe_dup_0[65]),.B2I1(NET_20),.B2I2(i_events[1]),.B2I3(NET_21),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.B2Z(NET_0),.Q2Z(i_events[1]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F13_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(i_events[4]),.T3I1(NET_20),.T3I2(fpgaio_oe_dup_0[68]),.T3I3(NET_21),.TB3S(GND),.C3Z(NET_667),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_F14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(lint_ADDR_int[3]),.B2I1(lint_ADDR_int[4]),.B2I2(NET_65),.B2I3(NET_68),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[3]),.T2I1(lint_ADDR_int[4]),.T2I2(NET_65),.T2I3(NET_68),.TB2S(lint_ADDR_int[6]),.C2Z(nx58292z1),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_F14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[66]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F15_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000010000000000),.B0I0(lint_ADDR_int[11]),.B0I1(NET_16),.B0I2(GND),.B0I3(NET_8),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.T0I0(NET_111),.T0I1(NET_129),.T0I2(fpgaio_in_int[28]),.T0I3(m1_m1_control[28]),.TB0S(GND),.B0Z(NET_128),.C0Z(NET_561),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F15_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[6]),.T1I1(NET_65),.T1I2(NET_67),.T1I3(NET_68),.C1Z(nx44608z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_F15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(m1_m1_sat_dup_0),.B2I1(fpgaio_in_int[18]),.B2I2(NET_111),.B2I3(NET_129),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.B2Z(NET_361),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F15_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_in_int[17]),.T3I1(m1_m1_clr_dup_0),.T3I2(NET_111),.T3I3(NET_129),.C3Z(NET_343),.Q3Z(m1_m1_control[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_F16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_128),.B0I1(m1_m1_tc_dup_0),.B0I2(NET_129),.B0I3(fpgaio_out_dup_0[70]),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.T0I0(NET_128),.T0I1(m1_m1_tc_dup_0),.T0I2(NET_129),.T0I3(fpgaio_out_dup_0[70]),.TB0S(NET_644),.C0Z(NET_641),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_340),.B1I1(NET_341),.B1I2(NET_343),.B1I3(NET_342),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.T1I0(NET_343),.T1I1(NET_342),.T1I2(NET_340),.T1I3(NET_341),.TB1S(NET_344),.C1Z(NET_331),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_F16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m1_m1_control[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_360),.B3I1(NET_361),.B3I2(NET_359),.B3I3(NET_358),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(NET_359),.T3I1(NET_358),.T3I2(NET_360),.T3I3(NET_361),.TB3S(NET_362),.C3Z(NET_350),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_F17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000001000000),.B0I0(GND),.B0I1(NET_31),.B0I2(NET_10),.B0I3(lint_ADDR_int[11]),.B0Z(NET_129),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_578),.B1I1(NET_577),.B1I2(NET_579),.B1I3(NET_576),.T1I0(NET_579),.T1I1(NET_576),.T1I2(NET_578),.T1I3(NET_577),.TB1S(NET_580),.C1Z(NET_568),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_F17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(fpgaio_out_dup_0[76]),.B2I1(m1_m1_mode_dup_0[0]),.B2I2(NET_129),.B2I3(NET_128),.T2I0(fpgaio_out_dup_0[76]),.T2I1(m1_m1_mode_dup_0[0]),.T2I2(NET_129),.T2I3(NET_128),.TB2S(NET_232),.C2Z(NET_229),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_F17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_561),.B3I1(NET_560),.B3I2(NET_558),.B3I3(NET_559),.T3I0(NET_558),.T3I1(NET_559),.T3I2(NET_561),.T3I3(NET_560),.TB3S(NET_562),.C3Z(NET_550),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_F18_0 (.tFragBitInfo(16'b0000000001101010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_3__CAND3_BLSTL_6_padClk),.QRT(not_RESET_3),.QST(GND),.T0I0(cnt3[2]),.T0I1(cnt3[0]),.T0I2(cnt3[1]),.T0I3(GND),.TB0S(GND),.Q0Z(cnt3[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_431),.B1I1(NET_432),.B1I2(NET_433),.B1I3(NET_434),.QCK(CLK_int_3__CAND3_BLSTL_6_padClk),.QRT(not_RESET_3),.QST(GND),.T1I0(NET_433),.T1I1(NET_434),.T1I2(NET_431),.T1I3(NET_432),.TB1S(NET_435),.C1Z(NET_423),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_F18_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_3__CAND3_BLSTL_6_padClk),.QRT(not_RESET_3),.QST(GND),.T2I0(GND),.T2I1(cnt3[0]),.T2I2(GND),.T2I3(GND),.TB2S(GND),.Q2Z(cnt3[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F18_3 (.tFragBitInfo(16'b0000000000010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_3__CAND3_BLSTL_6_padClk),.QRT(not_RESET_3),.QST(GND),.T3I0(GND),.T3I1(cnt3[0]),.T3I2(cnt3[1]),.T3I3(GND),.TB3S(GND),.Q3Z(cnt3[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F19_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_97),.B0I1(i_events[7]),.B0I2(fpgaio_out_dup_0[39]),.B0I3(NET_96),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T0I0(NET_97),.T0I1(fpgaio_out_dup_0[32]),.T0I2(i_events[0]),.T0I3(NET_96),.TB0S(GND),.B0Z(NET_466),.C0Z(NET_93),.Q0Z(i_events[7]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F19_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[6]),.T1I1(GND),.T1I2(lint_ADDR_int[5]),.T1I3(lint_ADDR_int[4]),.TB1S(GND),.C1Z(NET_98),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_F19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000000000000),.B2I0(lint_ADDR_int[11]),.B2I1(lint_ADDR_int[3]),.B2I2(NET_10),.B2I3(NET_98),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B2Z(NET_97),.Q2Z(i_events[0]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F19_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_out_dup_0[44]),.T3I1(NET_97),.T3I2(NET_96),.T3I3(i_events[12]),.C3Z(NET_220),.Q3Z(i_events[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_F20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_control[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F20_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_in_int[58]),.T1I1(NET_127),.T1I2(NET_119),.T1I3(m1_m0_control[26]),.C1Z(NET_527),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_F20_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[60]),.T2I1(NET_127),.T2I2(NET_119),.T2I3(m1_m0_control[28]),.TB2S(GND),.C2Z(NET_562),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_F20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(m1_m0_control[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(GND),.B0I1(lint_ADDR_int[19]),.B0I2(lint_ADDR_int[17]),.B0I3(lint_ADDR_int[18]),.B0Z(NET_143),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F21_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int[19]),.T3I1(lint_ADDR_int[16]),.T3I2(lint_ADDR_int[17]),.T3I3(lint_ADDR_int[18]),.C3Z(NET_73),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_F22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx4939z1_CAND4_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[39]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx4939z1_CAND4_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[63]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx4939z1_CAND4_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[51]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx4939z1_CAND4_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[46]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx4939z1_CAND4_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[40]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_127),.B0I1(m1_m0_sat_dup_0),.B0I2(NET_119),.B0I3(fpgaio_in_int[50]),.B0Z(NET_362),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F25_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_127),.T1I1(fpgaio_in_int[49]),.T1I2(NET_119),.T1I3(m1_m0_clr_dup_0),.C1Z(NET_344),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_F25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_clr_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_wdata_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_wdata_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[5]),.Q2EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_waddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wdata_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[11]),.Q0EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_waddr_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[6]),.Q1EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_waddr_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdata_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[4]),.Q3EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_waddr_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[7]),.Q0EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_waddr_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[3]),.Q1EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_waddr_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[1]),.Q2EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_waddr_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_waddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[9]),.Q0EN(nx34850z1_CAND5_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_raddr_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[0]),.Q1EN(nx34006z2_CAND2_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_waddr_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[10]),.Q2EN(nx34850z1_CAND5_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_raddr_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[6]),.Q3EN(nx34850z1_CAND5_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_raddr_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[11]),.Q0EN(nx34850z1_CAND5_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_raddr_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[11]),.Q1EN(nx34006z2_CAND2_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_waddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[7]),.Q2EN(nx34850z1_CAND5_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_raddr_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[8]),.Q3EN(nx34850z1_CAND5_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_raddr_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(NET_762),.Q2EN(nx34006z2_CAND2_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_we_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G5_0 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0000000000000000),.T0I0(lint_ADDR_int[12]),.T0I1(lint_ADDR_int[13]),.T0I2(NET_65),.T0I3(NET_144),.TB0S(GND),.C0Z(nx34006z2),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_G5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx39840z1_CAND4_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx39840z1_CAND4_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx39840z1_CAND4_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx39840z1_CAND4_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[19]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[73]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[78]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G12_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_20),.B0I1(i_events[11]),.B0I2(NET_21),.B0I3(fpgaio_oe_dup_0[75]),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.T0I0(NET_21),.T0I1(NET_20),.T0I2(fpgaio_oe_dup_0[67]),.T0I3(i_events[3]),.TB0S(GND),.B0Z(NET_193),.C0Z(NET_686),.Q0Z(i_events[11]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G12_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(NET_21),.T1I1(NET_20),.T1I2(i_events[13]),.T1I3(fpgaio_oe_dup_0[77]),.C1Z(NET_233),.Q1Z(i_events[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(i_events[14]),.B2I1(fpgaio_oe_dup_0[78]),.B2I2(NET_21),.B2I3(NET_20),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.B2Z(NET_253),.Q2Z(i_events[14]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.Q3Z(i_events[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G13_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.T0I0(RESET_int[2]),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND),.C0Z(not_RESET_2),.Q0Z(i_events[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G13_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(i_events[15]),.T1I1(NET_20),.T1I2(NET_21),.T1I3(fpgaio_oe_dup_0[79]),.TB1S(GND),.C1Z(NET_292),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_G13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000010000000),.B2I0(lint_ADDR_int[6]),.B2I1(lint_ADDR_int[3]),.B2I2(lint_ADDR_int[5]),.B2I3(lint_ADDR_int[4]),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.B2Z(NET_22),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G13_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(NET_22),.T3I1(NET_10),.T3I2(GND),.T3I3(GND),.C3Z(NET_21),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_5__CAND5_TLSBL_7_padClk),.QRT(not_RESET_2),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G14_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_5__CAND5_TLSBL_7_padClk),.QRT(not_RESET_2),.QST(GND),.T1I0(GND),.T1I1(GND),.T1I2(cnt5[0]),.T1I3(GND),.TB1S(GND),.Q1Z(cnt5[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_G14_2 (.tFragBitInfo(16'b0000000000010010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_5__CAND5_TLSBL_7_padClk),.QRT(not_RESET_2),.QST(GND),.T2I0(cnt5[1]),.T2I1(GND),.T2I2(cnt5[0]),.T2I3(GND),.TB2S(GND),.Q2Z(cnt5[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_G14_3 (.tFragBitInfo(16'b0001001100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_5__CAND5_TLSBL_7_padClk),.QRT(not_RESET_2),.QST(GND),.T3I0(cnt5[1]),.T3I1(GND),.T3I2(cnt5[0]),.T3I3(cnt5[2]),.TB3S(GND),.Q3Z(cnt5[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_G15_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_119),.B0I1(NET_118),.B0I2(m1_m0_outsel_dup_0[0]),.B0I3(fpgaio_in_int[64]),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.T0I0(NET_119),.T0I1(NET_118),.T0I2(m1_m0_mode_dup_0[0]),.T0I3(fpgaio_in_int[76]),.TB0S(GND),.B0Z(NET_104),.C0Z(NET_221),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G15_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(NET_102),.T1I1(m0_oper0_wmode_dup_0[0]),.T1I2(NET_103),.T1I3(fpgaio_out_dup_0[2]),.TB1S(GND),.C1Z(NET_710),.Q1Z(m0_m0_control[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_G15_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_102),.B2I1(fpgaio_out_dup_0[0]),.B2I2(NET_103),.B2I3(m0_oper0_rmode_dup_0[0]),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.T2I0(NET_119),.T2I1(NET_118),.T2I2(m1_m0_control[7]),.T2I3(fpgaio_in_int[71]),.TB2S(GND),.B2Z(NET_90),.C2Z(NET_467),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_G15_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(NET_102),.T3I1(m0_oper0_wdsel_dup_0),.T3I2(NET_103),.T3I3(fpgaio_out_dup_0[12]),.C3Z(NET_217),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G16_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_92),.B0I1(NET_93),.B0I2(NET_90),.B0I3(NET_91),.T0I0(NET_118),.T0I1(fpgaio_in_int[70]),.T0I2(m1_m0_tc_dup_0),.T0I3(NET_119),.TB0S(GND),.B0Z(NET_81),.C0Z(NET_633),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_G16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_379),.B1I1(NET_378),.B1I2(NET_377),.B1I3(NET_380),.T1I0(NET_377),.T1I1(NET_380),.T1I2(NET_379),.T1I3(NET_378),.TB1S(NET_381),.C1Z(NET_369),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_G16_2 (.tFragBitInfo(16'b0101010111111111),.bFragBitInfo(16'b0100010111001111),.B2I0(NET_94),.B2I1(lint_ADDR_int[11]),.B2I2(fpgaio_oe_dup_0[64]),.B2I3(m1_m0_dataout_int[0]),.T2I0(NET_94),.T2I1(lint_ADDR_int[11]),.T2I2(fpgaio_oe_dup_0[64]),.T2I3(m1_m0_dataout_int[0]),.TB2S(NET_20),.C2Z(NET_92),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_G16_3 (.tFragBitInfo(16'b0101010111111111),.bFragBitInfo(16'b0011111100010101),.B3I0(fpgaio_oe_dup_0[76]),.B3I1(m1_m0_dataout_int[12]),.B3I2(NET_94),.B3I3(lint_ADDR_int[11]),.T3I0(NET_94),.T3I1(lint_ADDR_int[11]),.T3I2(fpgaio_oe_dup_0[76]),.T3I3(m1_m0_dataout_int[12]),.TB3S(NET_20),.C3Z(NET_219),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_G17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_118),.B0I1(NET_108),.B0I2(cnt5[0]),.B0I3(m0_m0_control[28]),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T0I0(NET_118),.T0I1(NET_108),.T0I2(cnt5[0]),.T0I3(m0_m0_control[28]),.TB0S(NET_563),.C0Z(NET_559),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G17_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(NET_220),.T1I1(NET_217),.T1I2(NET_218),.T1I3(NET_219),.TB1S(GND),.C1Z(NET_215),.Q1Z(m0_m0_control[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_G17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_118),.B2I1(cnt5[1]),.B2I2(m0_m0_control[29]),.B2I3(NET_108),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(NET_118),.T2I1(cnt5[1]),.T2I2(m0_m0_control[29]),.T2I3(NET_108),.TB2S(NET_581),.C2Z(NET_577),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_G17_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_outsel_dup_0[2]),.T3I1(NET_118),.T3I2(fpgaio_in_int[66]),.T3I3(NET_119),.TB3S(GND),.C3Z(NET_714),.Q3Z(m0_m0_control[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_G18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(cnt3[1]),.B0I1(NET_108),.B0I2(m0_m0_control[23]),.B0I3(NET_118),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T0I0(cnt3[1]),.T0I1(NET_108),.T0I2(m0_m0_control[23]),.T0I3(NET_118),.TB0S(NET_454),.C0Z(NET_450),.Q0Z(m0_m0_control[24]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(cnt3[2]),.B1I1(NET_118),.B1I2(m0_m0_control[24]),.B1I3(NET_108),.CD1S(VCC),.Q1DI(lint_WDATA_int[23]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(m0_m0_control[24]),.T1I1(NET_108),.T1I2(cnt3[2]),.T1I3(NET_118),.TB1S(NET_493),.C1Z(NET_489),.Q1Z(m0_m0_control[23]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_G18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(cnt3[0]),.B2I1(NET_108),.B2I2(m0_m0_control[22]),.B2I3(NET_118),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(cnt3[0]),.T2I1(NET_108),.T2I2(m0_m0_control[22]),.T2I3(NET_118),.TB2S(NET_436),.C2Z(NET_432),.Q2Z(m0_oper0_wdsel_dup_0),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_G18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_control[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G19_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000010000000000),.B0I0(lint_ADDR_int[11]),.B0I1(NET_8),.B0I2(GND),.B0I3(NET_31),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_out_dup_0[34]),.T0I1(i_events[2]),.T0I2(NET_97),.T0I3(NET_96),.TB0S(GND),.B0Z(NET_119),.C0Z(NET_713),.Q0Z(i_events[2]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G19_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[38]),.T1I1(NET_96),.T1I2(NET_97),.T1I3(i_events[6]),.TB1S(GND),.C1Z(NET_632),.Q1Z(i_events[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_G19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx4939z1_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[56]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(m1_m0_control[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(m1_m1_control[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx4939z1_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[54]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G20_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(m1_m1_control[4]),.T2I1(NET_28),.T2I2(fpgaio_oe_dup_0[36]),.T2I3(NET_29_CAND5_BLSTL_7_tpGCLKBUF),.TB2S(GND),.C2Z(NET_674),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_G20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx4939z1_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[33]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_m1_control[10]),.B2I1(NET_29_CAND5_BLSTL_7_tpGCLKBUF),.B2I2(NET_28),.B2I3(fpgaio_oe_dup_0[42]),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B2Z(NET_181),.Q2Z(m1_m1_control[10]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wmode_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_rmode_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G22_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(NET_28),.T1I1(m1_m1_control[9]),.T1I2(fpgaio_oe_dup_0[41]),.T1I3(NET_29_CAND5_BLSTL_7_tpGCLKBUF),.C1Z(NET_159),.Q1Z(m1_m1_control[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_29_CAND5_BLSTL_7_tpGCLKBUF),.B2I1(fpgaio_oe_dup_0[37]),.B2I2(NET_28),.B2I3(m1_m1_control[5]),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B2Z(NET_654),.Q2Z(m1_m1_control[9]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx4939z1_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[59]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx4939z1_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[34]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx4939z1_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[38]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001000000000000),.B2I0(GND),.B2I1(lint_ADDR_int[13]),.B2I2(NET_65),.B2I3(NET_171),.B2Z(nx22245z1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_outsel_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(NET_762),.Q3EN(nx22245z1_CAND4_BLSBL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_we_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[6]),.Q0EN(nx60831z1_CAND3_BLSBL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_raddr_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[11]),.Q1EN(nx60831z1_CAND3_BLSBL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_raddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[5]),.Q2EN(nx60831z1_CAND3_BLSBL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_raddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[8]),.Q3EN(nx60831z1_CAND3_BLSBL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_raddr_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[7]),.Q0EN(nx60831z1_CAND3_BLSBL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_raddr_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[9]),.Q1EN(nx60831z1_CAND3_BLSBL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_raddr_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[10]),.Q2EN(nx60831z1_CAND3_BLSBL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_raddr_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[0]),.Q3EN(nx22245z1_CAND4_BLSBL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_waddr_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[4]),.Q0EN(nx34850z1_CAND5_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_raddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[1]),.Q1EN(nx34850z1_CAND5_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_raddr_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[5]),.Q2EN(nx34850z1_CAND5_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_raddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[0]),.Q3EN(nx34850z1_CAND5_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_raddr_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[3]),.Q0EN(nx34850z1_CAND5_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper0_raddr_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[2]),.Q2EN(nx34850z1_CAND5_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_raddr_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H5_0 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'b0000100000000000),.B0I0(NET_367),.B0I1(NET_142),.B0I2(GND),.B0I3(NET_141),.T0I0(lint_ADDR_int[13]),.T0I1(lint_ADDR_int[12]),.T0I2(lint_ADDR_int[14]),.T0I3(lint_WEN_int),.TB0S(GND),.B0Z(nx34850z1),.C0Z(NET_367),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_H5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx39840z1_CAND4_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[13]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H7_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_out_dup_0[3]),.T0I1(NET_61),.T0I2(m0_oper0_wmode_dup_0[1]),.T0I3(NET_60),.TB0S(GND),.C0Z(NET_703),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx39840z1_CAND4_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H7_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(NET_61),.T3I1(m0_oper0_rmode_dup_0[1]),.T3I2(fpgaio_out_dup_0[1]),.T3I3(NET_60),.C3Z(NET_56),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx39840z1_CAND4_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.QST(GND),.Q0Z(m0_m0_osel_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.QST(GND),.Q2Z(m0_m0_clr_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H11_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.QST(GND),.T0I0(m0_m0_outsel_dup_0[5]),.T0I1(NET_36),.T0I2(NET_37),.T0I3(fpgaio_in_int[69]),.TB0S(GND),.C0Z(NET_652),.Q0Z(m0_m0_sat_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H11_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_37),.T1I1(NET_36),.T1I2(fpgaio_in_int[73]),.T1I3(m0_m0_control[9]),.C1Z(NET_157),.Q1Z(m0_m0_control[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_H11_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.QST(GND),.T2I0(m0_m0_outsel_dup_0[3]),.T2I1(NET_36),.T2I2(NET_37),.T2I3(fpgaio_in_int[67]),.TB2S(GND),.C2Z(NET_691),.Q2Z(m0_m0_rnd_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_H11_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_in_int[75]),.T3I1(NET_36),.T3I2(NET_37),.T3I3(m0_m0_control[11]),.TB3S(GND),.C3Z(NET_198),.Q3Z(m0_m0_control[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_H12_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_36),.B0I1(fpgaio_in_int[78]),.B0I2(m0_m0_osel_dup_0),.B0I3(NET_37),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_4__CAND4_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T0I0(GND),.T0I1(cnt4[0]),.T0I2(GND),.T0I3(GND),.TB0S(GND),.B0Z(NET_258),.Q0Z(cnt4[0]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H12_1 (.tFragBitInfo(16'b0001010101000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_4__CAND4_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T1I0(GND),.T1I1(cnt4[0]),.T1I2(cnt4[1]),.T1I3(cnt4[2]),.TB1S(GND),.Q1Z(cnt4[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H12_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_37),.B2I1(cnt4[0]),.B2I2(fpgaio_out_dup_0[25]),.B2I3(NET_60),.QCK(CLK_int_4__CAND4_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T2I0(cnt2[1]),.T2I1(NET_37),.T2I2(fpgaio_out_dup_0[20]),.T2I3(NET_60),.TB2S(GND),.B2Z(NET_510),.C2Z(NET_400),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_H12_3 (.tFragBitInfo(16'b0000000000010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_4__CAND4_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T3I0(GND),.T3I1(cnt4[0]),.T3I2(cnt4[1]),.T3I3(GND),.TB3S(GND),.Q3Z(cnt4[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_H13_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001000000000000),.B0I0(GND),.B0I1(GND),.B0I2(NET_22),.B0I3(NET_8),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T0I0(cnt5[2]),.T0I1(NET_60),.T0I2(fpgaio_out_dup_0[30]),.T0I3(NET_37),.TB0S(GND),.B0Z(NET_37),.C0Z(NET_598),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H13_1 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T1I0(lint_ADDR_int[5]),.T1I1(lint_ADDR_int[3]),.T1I2(lint_ADDR_int[4]),.T1I3(lint_ADDR_int[6]),.C1Z(NET_16),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_H13_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T2I0(cnt1[0]),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND),.Q2Z(cnt1[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_H13_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T3I0(cnt1[0]),.T3I1(NET_60),.T3I2(fpgaio_out_dup_0[16]),.T3I3(NET_37),.TB3S(GND),.C3Z(NET_326),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_H14_0 (.tFragBitInfo(16'b0000000001101100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T0I0(cnt1[0]),.T0I1(cnt1[2]),.T0I2(cnt1[1]),.T0I3(GND),.TB0S(GND),.Q0Z(cnt1[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(NET_118),.B1I1(cnt1[2]),.B1I2(NET_108),.B1I3(m0_m0_sat_dup_0),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T1I0(NET_108),.T1I1(m0_m0_sat_dup_0),.T1I2(NET_118),.T1I3(cnt1[2]),.TB1S(NET_363),.C1Z(NET_359),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_H14_2 (.tFragBitInfo(16'b0000000000000110),.bFragBitInfo(16'b0000001000000000),.B2I0(NET_22),.B2I1(lint_ADDR_int[11]),.B2I2(GND),.B2I3(NET_8),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T2I0(cnt1[0]),.T2I1(cnt1[1]),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(NET_118),.Q2Z(cnt1[1]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_H14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B3I0(NET_118),.B3I1(m0_m0_clr_dup_0),.B3I2(NET_108),.B3I3(cnt1[1]),.QCK(CLK_int_1__CAND1_TLSBL_8_padClk),.QRT(not_RESET_1),.QST(GND),.T3I0(NET_108),.T3I1(cnt1[1]),.T3I2(NET_118),.T3I3(m0_m0_clr_dup_0),.TB3S(NET_345),.C3Z(NET_341),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_H15_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000011101110111),.B0I0(m0_oper1_wmode_dup_0[1]),.B0I1(NET_103),.B0I2(fpgaio_out_dup_0[7]),.B0I3(NET_102),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_2__CAND2_TLSBL_8_padClk),.QRT(not_RESET_2),.QST(GND),.T0I0(GND),.T0I1(cnt2[0]),.T0I2(GND),.T0I3(GND),.TB0S(GND),.B0Z(NET_463),.Q0Z(cnt2[0]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H15_1 (.tFragBitInfo(16'b0001010101000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_2__CAND2_TLSBL_8_padClk),.QRT(not_RESET_2),.QST(GND),.T1I0(GND),.T1I1(cnt2[0]),.T1I2(cnt2[1]),.T1I3(cnt2[2]),.TB1S(GND),.Q1Z(cnt2[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_108),.B2I1(cnt2[0]),.B2I2(m0_m0_control[19]),.B2I3(NET_118),.QCK(CLK_int_2__CAND2_TLSBL_8_padClk),.QRT(not_RESET_2),.QST(GND),.T2I0(NET_108),.T2I1(cnt2[0]),.T2I2(m0_m0_control[19]),.T2I3(NET_118),.TB2S(NET_382),.C2Z(NET_378),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_H15_3 (.tFragBitInfo(16'b0000000000010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_2__CAND2_TLSBL_8_padClk),.QRT(not_RESET_2),.QST(GND),.T3I0(GND),.T3I1(cnt2[0]),.T3I2(cnt2[1]),.T3I3(GND),.TB3S(GND),.Q3Z(cnt2[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_H16_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.T0I0(NET_80),.T0I1(NET_81),.T0I2(NET_78),.T0I3(NET_79),.TB0S(GND),.Q0Z(lint_RDATA_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H16_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.T1I0(NET_466),.T1I1(NET_463),.T1I2(NET_465),.T1I3(NET_464),.TB1S(GND),.C1Z(NET_461),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_H16_2 (.tFragBitInfo(16'b0101111101011111),.bFragBitInfo(16'b0101111100010011),.B2I0(NET_94),.B2I1(fpgaio_oe_dup_0[71]),.B2I2(m1_m0_dataout_int[7]),.B2I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.T2I0(NET_94),.T2I1(fpgaio_oe_dup_0[71]),.T2I2(m1_m0_dataout_int[7]),.T2I3(lint_ADDR_int[11]),.TB2S(NET_20),.C2Z(NET_465),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_H16_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF),.T3I0(NET_460),.T3I1(NET_458),.T3I2(NET_461),.T3I3(NET_459),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_H17_0 (.tFragBitInfo(16'b0011001111111111),.bFragBitInfo(16'b0010001110101111),.B0I0(lint_ADDR_int[11]),.B0I1(m1_m0_dataout_int[2]),.B0I2(fpgaio_oe_dup_0[66]),.B0I3(NET_94),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.T0I0(lint_ADDR_int[11]),.T0I1(m1_m0_dataout_int[2]),.T0I2(fpgaio_oe_dup_0[66]),.T0I3(NET_94),.TB0S(NET_20),.C0Z(NET_712),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H17_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.T1I0(NET_712),.T1I1(NET_713),.T1I2(NET_711),.T1I3(NET_710),.C1Z(NET_708),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_H17_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.T2I0(NET_707),.T2I1(NET_706),.T2I2(NET_708),.T2I3(NET_705),.TB2S(GND),.Q2Z(lint_RDATA_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_H17_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.T3I0(NET_214),.T3I1(NET_212),.T3I2(NET_215),.T3I3(NET_213),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_H18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q0Z(m0_m0_control[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_524),.B1I1(NET_526),.B1I2(NET_525),.B1I3(NET_523),.CD1S(VCC),.Q1DI(lint_WDATA_int[26]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_525),.T1I1(NET_523),.T1I2(NET_524),.T1I3(NET_526),.TB1S(NET_527),.C1Z(NET_515),.Q1Z(m0_m0_control[26]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_H18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(cnt4[1]),.B2I1(NET_108),.B2I2(NET_118),.B2I3(m0_m0_control[26]),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T2I0(cnt4[1]),.T2I1(NET_108),.T2I2(NET_118),.T2I3(m0_m0_control[26]),.TB2S(NET_528),.C2Z(NET_524),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_H18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(NET_118),.B3I1(NET_108),.B3I2(cnt2[2]),.B3I3(m0_m0_control[21]),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(cnt2[2]),.T3I1(m0_m0_control[21]),.T3I2(NET_118),.T3I3(NET_108),.TB3S(NET_418),.C3Z(NET_414),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_H19_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(apb_fsm[1]),.TB0S(GND),.C0Z(not_apb_fsm_1),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_rmode_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000100),.B2I0(lint_GNT_dup_0),.B2I1(lint_REQ_int),.B2I2(apb_fsm[0]),.B2I3(apb_fsm[1]),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B2Z(NET_142),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H19_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx4939z1_CAND4_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[2]),.T3I1(lint_ADDR_int[6]),.T3I2(NET_65),.T3I3(GND),.TB3S(GND),.C3Z(NET_602),.Q3Z(fpgaio_out_dup_0[47]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_H20_0 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx4939z1_CAND4_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(lint_WEN_int),.T0I1(GND),.T0I2(lint_GNT_dup_0),.T0I3(lint_REQ_int),.TB0S(GND),.C0Z(nx7012z2),.Q0Z(fpgaio_out_dup_0[45]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H20_1 (.tFragBitInfo(16'b1110111111101110),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T1I0(apb_fsm[0]),.T1I1(apb_fsm[1]),.T1I2(lint_GNT_dup_0),.T1I3(lint_REQ_int),.TB1S(GND),.C1Z(nx10146z2),.Q1Z(m0_oper0_wmode_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_H20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001001),.B2I0(apb_fsm[0]),.B2I1(apb_fsm[1]),.B2I2(GND),.B2I3(GND),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B2Z(nx7012z3),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H20_3 (.tFragBitInfo(16'b0000000000001110),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3EN(nx7012z3),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(nx7012z2),.T3I1(apb_fsm[1]),.T3I2(GND),.T3I3(GND),.TB3S(GND),.Q3Z(lint_GNT_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.Q3DI(GND),.T3CO());

	LOGIC_0 QL_INST_H21_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000001000),.B0I0(lint_ADDR_int[12]),.B0I1(lint_ADDR_int[14]),.B0I2(lint_ADDR_int[15]),.B0I3(lint_ADDR_int[16]),.CD0S(VCC),.Q0DI(lint_WDATA_int[28]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(m1_m0_dataout_int[29]),.T0I1(NET_94),.T0I2(m0_ram_control[29]),.T0I3(NET_103),.TB0S(GND),.B0Z(NET_252),.C0Z(NET_573),.Q0Z(m0_ram_control[28]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx4939z1_CAND4_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[48]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H21_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000010000),.B2I0(lint_ADDR_int[15]),.B2I1(lint_ADDR_int[14]),.B2I2(NET_143),.B2I3(lint_ADDR_int[16]),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T2I0(m1_m0_dataout_int[28]),.T2I1(m0_ram_control[28]),.T2I2(NET_94),.T2I3(NET_103),.TB2S(GND),.B2Z(NET_144),.C2Z(NET_555),.Q2Z(m0_ram_control[29]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_H21_3 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[15]),.T3I1(GND),.T3I2(NET_143),.T3I3(lint_ADDR_int[16]),.C3Z(NET_141),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_29_CAND5_BLSTL_8_tpGCLKBUF),.B0I1(NET_28),.B0I2(fpgaio_oe_dup_0[43]),.B0I3(m1_m1_control[11]),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0Z(NET_200),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_control[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_outsel_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H23_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_WEN_int),.T1I1(lint_ADDR_int[13]),.T1I2(NET_171),.T1I3(NET_142),.TB1S(GND),.C1Z(nx60831z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_H23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx4939z1_CAND4_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[60]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx4939z1_CAND4_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[61]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[18]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_sat_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_rnd_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_outsel_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_osel_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[4]),.Q1EN(nx60831z1_CAND3_BLSBL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_raddr_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[2]),.Q2EN(nx60831z1_CAND3_BLSBL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_raddr_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[3]),.Q0EN(nx60831z1_CAND3_BLSBL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper0_raddr_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[0]),.Q1EN(nx60831z1_CAND3_BLSBL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper0_raddr_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[1]),.Q3EN(nx60831z1_CAND3_BLSBL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_raddr_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I3_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_oe_dup_0[9]),.B0I1(m0_m0_dataout_int[9]),.B0I2(NET_58),.B0I3(NET_59),.T0I0(fpgaio_oe_dup_0[1]),.T0I1(m0_m0_dataout_int[1]),.T0I2(NET_58),.T0I3(NET_59),.TB0S(GND),.B0Z(NET_168),.C0Z(NET_55),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_I3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I3_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_59),.T3I1(fpgaio_oe_dup_0[3]),.T3I2(NET_58),.T3I3(m0_m0_dataout_int[3]),.TB3S(GND),.C3Z(NET_702),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_I7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_54),.B0I1(NET_55),.B0I2(NET_53),.B0I3(NET_56),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND3_TLSTR_9_tpGCLKBUF),.QST(GND),.B0Z(NET_57),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I7_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND3_TLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_701),.T1I1(NET_700),.T1I2(NET_703),.T1I3(NET_702),.TB1S(GND),.C1Z(NET_704),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_I7_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND3_TLSTR_9_tpGCLKBUF),.QST(GND),.T2I0(m0_coef_rmode_dup_0[1]),.T2I1(NET_60),.T2I2(fpgaio_out_dup_0[9]),.T2I3(NET_61),.TB2S(GND),.C2Z(NET_169),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I7_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND3_TLSTR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_168),.T3I1(NET_169),.T3I2(NET_167),.T3I3(NET_166),.TB3S(GND),.C3Z(NET_170),.Q3Z(fpgaio_out_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_I10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[65]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.Q2Z(m0_m0_outsel_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[67]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I11_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000001),.B0I0(lint_ADDR_int[7]),.B0I1(lint_ADDR_int[8]),.B0I2(apb_fsm[0]),.B0I3(lint_ADDR_int[2]),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T0I0(m0_m0_outsel_dup_0[1]),.T0I1(NET_37),.T0I2(fpgaio_in_int[65]),.T0I3(NET_36),.TB0S(GND),.B0Z(NET_8),.C0Z(NET_23),.Q0Z(m0_m0_control[8]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[79]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I11_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(NET_36),.T2I1(NET_37),.T2I2(fpgaio_in_int[68]),.T2I3(m0_m0_outsel_dup_0[4]),.TB2S(GND),.C2Z(NET_672),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I11_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_control[8]),.T3I1(NET_37),.T3I2(fpgaio_in_int[72]),.T3I3(NET_36),.TB3S(GND),.C3Z(NET_278),.Q3Z(fpgaio_out_dup_0[72]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_I12_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T0I0(cnt4[2]),.T0I1(NET_37),.T0I2(NET_60),.T0I3(fpgaio_out_dup_0[27]),.TB0S(GND),.C0Z(NET_545),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I12_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_36),.T1I1(NET_37),.T1I2(m0_m0_control[10]),.T1I3(fpgaio_in_int[74]),.TB1S(GND),.C1Z(NET_179),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_I12_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[77]),.T2I1(NET_36),.T2I2(NET_37),.T2I3(m0_m0_mode_dup_0[1]),.TB2S(GND),.C2Z(NET_238),.Q2Z(m0_m0_csel_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_I12_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_36),.T3I1(NET_37),.T3I2(m0_m0_csel_dup_0),.T3I3(fpgaio_in_int[79]),.TB3S(GND),.C3Z(NET_297),.Q3Z(m0_m0_control[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_I13_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(saved_REQ),.B0I1(fpgaio_out_dup_0[31]),.B0I2(NET_37),.B0I3(NET_60),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.T0I0(NET_692),.T0I1(NET_691),.T0I2(NET_694),.T0I3(NET_693),.TB0S(GND),.B0Z(NET_616),.C0Z(NET_695),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I13_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.T1I0(NET_160),.T1I1(NET_157),.T1I2(NET_158),.T1I3(NET_159),.TB1S(GND),.C1Z(NET_161),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_I13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I13_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_730),.B3I1(NET_161),.B3I2(NET_164),.B3I3(NET_156),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64_CAND2_TLSBR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.T3I0(NET_164),.T3I1(NET_156),.T3I2(NET_730),.T3I3(NET_161),.TB3S(NET_170),.Q3Z(lint_RDATA_dup_0[9]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_I14_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B0I0(fpgaio_out_dup_0[22]),.B0I1(NET_85),.B0I2(m1_ram_control[22]),.B0I3(NET_102),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T0I0(NET_85),.T0I1(fpgaio_out_dup_0[24]),.T0I2(m1_ram_control[24]),.T0I3(NET_102),.TB0S(GND),.B0Z(NET_429),.C0Z(NET_486),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I14_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_85),.T1I1(fpgaio_out_dup_0[26]),.T1I2(m1_ram_control[26]),.T1I3(NET_102),.TB1S(GND),.C1Z(NET_521),.Q1Z(m1_ram_control[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_I14_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[6]),.T2I1(NET_65),.T2I2(NET_68),.T2I3(NET_146),.TB2S(GND),.C2Z(nx39840z1),.Q2Z(m1_ram_control[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_I14_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_645),.T3I1(lint_ADDR_int[4]),.T3I2(NET_68),.T3I3(lint_ADDR_int[6]),.TB3S(GND),.C3Z(nx53524z1),.Q3Z(m1_ram_control[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_I15_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000010000000),.B0I0(NET_8),.B0I1(NET_11),.B0I2(NET_9),.B0I3(GND),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T0I0(m1_ram_control[29]),.T0I1(NET_102),.T0I2(fpgaio_out_dup_0[29]),.T0I3(NET_85),.TB0S(GND),.B0Z(NET_60),.C0Z(NET_574),.Q0Z(m1_ram_control[29]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I15_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[23]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[23]),.T1I1(NET_102),.T1I2(m1_ram_control[23]),.T1I3(NET_85),.TB1S(GND),.C1Z(NET_447),.Q1Z(m1_ram_control[23]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_I15_2 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_9),.B2I1(NET_8),.B2I2(GND),.B2I3(NET_88),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_ADDR_int[5]),.T2I2(GND),.T2I3(lint_ADDR_int[6]),.TB2S(GND),.B2Z(NET_102),.C2Z(NET_9),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I15_3 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_10),.T3I1(lint_ADDR_int[5]),.T3I2(lint_ADDR_int[6]),.T3I3(NET_88),.TB3S(GND),.C3Z(NET_85),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_I16_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000100000000000),.B0I0(NET_8),.B0I1(lint_ADDR_int[5]),.B0I2(lint_ADDR_int[6]),.B0I3(NET_88),.T0I0(GND),.T0I1(lint_ADDR_int[3]),.T0I2(lint_ADDR_int[11]),.T0I3(lint_ADDR_int[4]),.TB0S(GND),.B0Z(NET_103),.C0Z(NET_88),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_I16_1 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(GND),.T1I1(NET_88),.T1I2(NET_9),.T1I3(NET_10),.TB1S(GND),.C1Z(NET_96),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_I16_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_8),.B2I1(lint_ADDR_int[3]),.B2I2(NET_9),.B2I3(lint_ADDR_int[4]),.T2I0(NET_629),.T2I1(NET_632),.T2I2(NET_630),.T2I3(NET_631),.TB2S(GND),.B2Z(NET_20),.C2Z(NET_627),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_I16_3 (.tFragBitInfo(16'b0111011101110111),.bFragBitInfo(16'b0000101110111011),.B3I0(lint_ADDR_int[11]),.B3I1(fpgaio_oe_dup_0[70]),.B3I2(m1_m0_dataout_int[6]),.B3I3(NET_94),.T3I0(m1_m0_dataout_int[6]),.T3I1(NET_94),.T3I2(lint_ADDR_int[11]),.T3I3(fpgaio_oe_dup_0[70]),.TB3S(NET_20),.C3Z(NET_631),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_I17_0 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0100000000000000),.B0I0(GND),.B0I1(NET_9),.B0I2(NET_10),.B0I3(NET_11),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.T0I0(NET_519),.T0I1(GND),.T0I2(NET_521),.T0I3(NET_520),.TB0S(GND),.B0Z(NET_5),.C0Z(NET_517),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I17_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.T1I0(NET_573),.T1I1(GND),.T1I2(NET_574),.T1I3(NET_572),.TB1S(GND),.C1Z(NET_570),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_I17_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.T2I0(NET_569),.T2I1(NET_567),.T2I2(NET_568),.T2I3(NET_570),.TB2S(GND),.Q2Z(lint_RDATA_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_I17_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.T3I0(NET_517),.T3I1(NET_515),.T3I2(NET_516),.T3I3(NET_514),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_I18_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.T0I0(NET_441),.T0I1(NET_440),.T0I2(NET_442),.T0I3(NET_443),.TB0S(GND),.Q0Z(lint_RDATA_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I18_1 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.T1I0(GND),.T1I1(NET_445),.T1I2(NET_447),.T1I3(NET_446),.TB1S(GND),.C1Z(NET_443),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_I18_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0100000000000000),.B2I0(GND),.B2I1(NET_429),.B2I2(NET_427),.B2I3(NET_428),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.T2I0(NET_485),.T2I1(NET_486),.T2I2(GND),.T2I3(NET_484),.TB2S(GND),.B2Z(NET_425),.C2Z(NET_482),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I18_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.T3I0(NET_479),.T3I1(NET_480),.T3I2(NET_482),.T3I3(NET_481),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_I19_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(GND),.T0I0(GND),.T0I1(GND),.T0I2(lint_ADDR_int[4]),.T0I3(lint_ADDR_int[3]),.TB0S(GND),.C0Z(NET_11),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I19_1 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(GND),.T1I0(lint_ADDR_int[6]),.T1I1(lint_ADDR_int[5]),.T1I2(lint_ADDR_int[4]),.T1I3(lint_ADDR_int[3]),.TB1S(GND),.C1Z(NET_31),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_I19_2 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_REQ_int),.Q2EN(RESET_int[0]),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(GND),.T2I0(lint_ADDR_int[6]),.T2I1(lint_ADDR_int[5]),.T2I2(NET_8),.T2I3(NET_11),.TB2S(GND),.C2Z(NET_61),.Q2Z(saved_REQ),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_I19_3 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(GND),.QST(GND),.T3I0(NET_10),.T3I1(GND),.T3I2(NET_31),.T3I3(GND),.TB3S(GND),.C3Z(NET_28),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_I20_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_5),.B0I1(m0_m0_dataout_int[25]),.B0I2(NET_59),.B0I3(fpgaio_out_dup_0[57]),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T0I0(NET_5),.T0I1(fpgaio_out_dup_0[59]),.T0I2(NET_59),.T0I3(m0_m0_dataout_int[27]),.TB0S(GND),.B0Z(NET_502),.C0Z(NET_537),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I20_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(apb_fsm[0]),.T1I2(GND),.T1I3(GND),.C1Z(not_apb_fsm_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_I20_2 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'b0000000000000001),.B2I0(lint_WEN_int),.B2I1(apb_fsm[0]),.B2I2(GND),.B2I3(GND),.CD2S(GND),.Q2EN(nx10146z2),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T2I0(nx10146z1),.T2I1(GND),.T2I2(apb_fsm[1]),.T2I3(not_apb_fsm_0),.TB2S(GND),.B2Z(nx10146z1),.Q2Z(apb_fsm[0]),.B2CO(),.C2Z(),.Q2DI(GND),.T2CO());

	LOGIC_3 QL_INST_I20_3 (.tFragBitInfo(16'b0000000000110010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx10146z2),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T3I0(lint_WEN_int),.T3I1(apb_fsm[0]),.T3I2(apb_fsm[1]),.T3I3(GND),.TB3S(GND),.Q3Z(apb_fsm[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_I21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001000),.B0I0(lint_ADDR_int[14]),.B0I1(NET_73),.B0I2(lint_ADDR_int[12]),.B0I3(lint_ADDR_int[15]),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B0Z(NET_171),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I21_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[26]),.Q1EN(nx19726z1_CAND2_BLSTR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_59),.T1I1(fpgaio_out_dup_0[62]),.T1I2(NET_5),.T1I3(m0_m0_dataout_int[30]),.TB1S(GND),.C1Z(NET_590),.Q1Z(m0_ram_control[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_I21_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_m0_dataout_int[24]),.B2I1(NET_94),.B2I2(m0_ram_control[24]),.B2I3(NET_103),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T2I0(NET_59),.T2I1(NET_5),.T2I2(m0_m0_dataout_int[31]),.T2I3(fpgaio_out_dup_0[63]),.TB2S(GND),.B2Z(NET_485),.C2Z(NET_608),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I21_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[24]),.Q3EN(nx19726z1_CAND2_BLSTR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_94),.T3I1(m1_m0_dataout_int[26]),.T3I2(m0_ram_control[26]),.T3I3(NET_103),.C3Z(NET_520),.Q3Z(m0_ram_control[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_I22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[22]),.Q0EN(nx19726z1_CAND2_BLSTR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q0Z(m0_ram_control[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_control[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I22_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_94),.B2I1(NET_103),.B2I2(m0_ram_control[23]),.B2I3(m1_m0_dataout_int[23]),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T2I0(NET_28_CAND4_BLSTR_9_tpGCLKBUF),.T2I1(NET_29),.T2I2(fpgaio_oe_dup_0[35]),.T2I3(m1_m1_control[3]),.TB2S(GND),.B2Z(NET_446),.C2Z(NET_693),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I22_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx19726z1_CAND2_BLSTR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_94),.T3I1(m1_m0_dataout_int[22]),.T3I2(m0_ram_control[22]),.T3I3(NET_103),.TB3S(GND),.C3Z(NET_428),.Q3Z(m0_ram_control[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_I23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[42]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_mode_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_outsel_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J3_0 (.tFragBitInfo(16'b1111111101010101),.bFragBitInfo(16'b1111110001010101),.B0I0(lint_ADDR_int[11]),.B0I1(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.B0I2(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.B0I3(apb_fsm[0]),.T0I0(lint_ADDR_int[11]),.T0I1(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.T0I2(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.T0I3(apb_fsm[0]),.TB0S(m0_oper0_rdata_int[8]),.C0Z(NET_286),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J3_1 (.tFragBitInfo(16'b1111111101010101),.bFragBitInfo(16'b1100111110001011),.B1I0(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.B1I1(apb_fsm[0]),.B1I2(lint_ADDR_int[11]),.B1I3(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.T1I0(lint_ADDR_int[11]),.T1I1(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.T1I2(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.T1I3(apb_fsm[0]),.TB1S(m0_oper0_rdata_int[5]),.C1Z(NET_660),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_J3_2 (.tFragBitInfo(16'b1111111101010101),.bFragBitInfo(16'b1111110001010101),.B2I0(lint_ADDR_int[11]),.B2I1(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.B2I2(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.B2I3(apb_fsm[0]),.T2I0(lint_ADDR_int[11]),.T2I1(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.T2I2(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.T2I3(apb_fsm[0]),.TB2S(m0_oper0_rdata_int[9]),.C2Z(NET_165),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J3_3 (.tFragBitInfo(16'b1111111101010101),.bFragBitInfo(16'b1100111110001011),.B3I0(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.B3I1(apb_fsm[0]),.B3I2(lint_ADDR_int[11]),.B3I3(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.T3I0(lint_ADDR_int[11]),.T3I1(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.T3I2(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.T3I3(apb_fsm[0]),.TB3S(m0_oper0_rdata_int[13]),.C3Z(NET_246),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J4_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_58),.B0I1(fpgaio_oe_dup_0[14]),.B0I2(NET_59),.B0I3(m0_m0_dataout_int[14]),.T0I0(NET_58),.T0I1(m0_m0_dataout_int[15]),.T0I2(NET_59),.T0I3(fpgaio_oe_dup_0[15]),.TB0S(GND),.B0Z(NET_269),.C0Z(NET_308),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J4_1 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1110000011101111),.B1I0(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.B1I1(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.B1I2(apb_fsm[0]),.B1I3(lint_ADDR_int[11]),.T1I0(apb_fsm[0]),.T1I1(lint_ADDR_int[11]),.T1I2(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.T1I3(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.TB1S(m0_oper0_rdata_int[15]),.C1Z(NET_305),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_J4_2 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1011101110110001),.B2I0(apb_fsm[0]),.B2I1(lint_ADDR_int[11]),.B2I2(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.B2I3(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.T2I0(apb_fsm[0]),.T2I1(lint_ADDR_int[11]),.T2I2(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.T2I3(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.TB2S(m0_oper0_rdata_int[4]),.C2Z(NET_680),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J4_3 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1110000011101111),.B3I0(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.B3I1(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.B3I2(apb_fsm[0]),.B3I3(lint_ADDR_int[11]),.T3I0(apb_fsm[0]),.T3I1(lint_ADDR_int[11]),.T3I2(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.T3I3(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.TB3S(m0_oper0_rdata_int[11]),.C3Z(NET_206),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J5_2 (.tFragBitInfo(16'b1101110111011101),.bFragBitInfo(16'b1101110111010001),.B2I0(lint_ADDR_int[11]),.B2I1(apb_fsm[0]),.B2I2(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.B2I3(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.T2I0(lint_ADDR_int[11]),.T2I1(apb_fsm[0]),.T2I2(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF),.T2I3(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF),.TB2S(m0_oper0_rdata_int[3]),.C2Z(NET_699),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J7_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.T0I0(NET_267),.T0I1(NET_270),.T0I2(NET_268),.T0I3(NET_269),.TB0S(GND),.C0Z(NET_271),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_307),.B0I1(NET_308),.B0I2(NET_309),.B0I3(NET_306),.B0Z(NET_310),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(fpgaio_out_dup_0[15]),.B2I1(NET_61),.B2I2(m0_ram_control[15]),.B2I3(NET_60),.B2Z(NET_309),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J10_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.T0I0(fpgaio_out_dup_0[65]),.T0I1(tcdm_result_p0[1]),.T0I2(NET_12),.T0I3(NET_13),.TB0S(GND),.C0Z(NET_3),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J10_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(tcdm_result_p0[3]),.T3I1(NET_13),.T3I2(NET_12),.T3I3(fpgaio_out_dup_0[67]),.C3Z(NET_689),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J11_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_27),.B0I1(NET_728),.B0I2(NET_42),.B0I3(NET_4),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64_CAND2_TLSBR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T0I0(NET_27),.T0I1(NET_728),.T0I2(NET_42),.T0I3(NET_4),.TB0S(NET_57),.Q0Z(lint_RDATA_dup_0[1]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J11_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T1I0(NET_12),.T1I1(fpgaio_out_dup_0[79]),.T1I2(NET_13),.T1I3(tcdm_result_p0[15]),.TB1S(GND),.C1Z(NET_295),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_J11_2 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_12),.B2I1(fpgaio_out_dup_0[73]),.B2I2(NET_13),.B2I3(tcdm_result_p0[9]),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T2I0(NET_8),.T2I1(NET_16),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(NET_155),.C2Z(NET_12),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J11_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T3I0(NET_12),.T3I1(fpgaio_out_dup_0[78]),.T3I2(NET_13),.T3I3(tcdm_result_p0[14]),.C3Z(NET_256),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J12_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_265),.B0I1(NET_262),.B0I2(NET_257),.B0I3(NET_738),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64_CAND2_TLSBR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T0I0(NET_265),.T0I1(NET_262),.T0I2(NET_257),.T0I3(NET_738),.TB0S(NET_271),.Q0Z(lint_RDATA_dup_0[14]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J12_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B1I0(NET_690),.B1I1(NET_698),.B1I2(NET_761),.B1I3(NET_695),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64_CAND2_TLSBR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T1I0(NET_761),.T1I1(NET_695),.T1I2(NET_690),.T1I3(NET_698),.TB1S(NET_704),.Q1Z(lint_RDATA_dup_0[3]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_J12_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_256),.B2I1(NET_253),.B2I2(NET_255),.B2I3(NET_254),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T2I0(NET_689),.T2I1(NET_687),.T2I2(NET_686),.T2I3(NET_688),.TB2S(GND),.B2Z(NET_257),.C2Z(NET_690),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J13_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_154),.B0I1(NET_155),.B0I2(NET_153),.B0I3(NET_152),.T0I0(NET_36),.T0I1(NET_6),.T0I2(m0_m0_rnd_dup_0),.T0I3(tcdm_rdata_p2_int[16]),.TB0S(GND),.B0Z(NET_156),.C0Z(NET_329),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J13_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_2),.T1I1(NET_3),.T1I2(NET_0),.T1I3(NET_1),.C1Z(NET_4),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J13_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_328),.T2I1(NET_326),.T2I2(NET_327),.T2I3(NET_329),.TB2S(GND),.C2Z(NET_313),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J13_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_293),.T3I1(NET_294),.T3I2(NET_295),.T3I3(NET_292),.TB3S(GND),.C3Z(NET_296),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J14_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.QST(GND),.T0I0(NET_102),.T0I1(fpgaio_out_dup_0[19]),.T0I2(NET_85),.T0I3(m1_ram_control[19]),.TB0S(GND),.C0Z(NET_375),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J14_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_672),.T1I1(NET_675),.T1I2(NET_674),.T1I3(NET_673),.TB1S(GND),.C1Z(NET_676),.Q1Z(m1_ram_control[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_J14_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_23),.B2I1(NET_25),.B2I2(NET_24),.B2I3(NET_26),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.QST(GND),.T2I0(NET_261),.T2I1(NET_259),.T2I2(NET_260),.T2I3(NET_258),.TB2S(GND),.B2Z(NET_27),.C2Z(NET_262),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J14_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(RESET_int[1]),.T3I2(GND),.T3I3(GND),.TB3S(GND),.C3Z(not_RESET_1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_J15_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B0I0(m1_ram_control[28]),.B0I1(NET_85),.B0I2(NET_102),.B0I3(fpgaio_out_dup_0[28]),.CD0S(VCC),.Q0DI(lint_WDATA_int[28]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.QST(GND),.T0I0(NET_103),.T0I1(fpgaio_out_dup_0[6]),.T0I2(NET_102),.T0I3(m0_oper1_wmode_dup_0[0]),.TB0S(GND),.B0Z(NET_556),.C0Z(NET_629),.Q0Z(m1_ram_control[28]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J15_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[21]),.T1I1(NET_85),.T1I2(NET_102),.T1I3(m1_ram_control[21]),.TB1S(GND),.C1Z(NET_411),.Q1Z(m1_ram_control[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_J15_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.QST(GND),.T2I0(m1_ram_control[17]),.T2I1(fpgaio_out_dup_0[17]),.T2I2(NET_102),.T2I3(NET_85),.TB2S(GND),.C2Z(NET_338),.Q2Z(m1_ram_control[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_J15_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_out_dup_0[18]),.T3I1(NET_85),.T3I2(NET_102),.T3I3(m1_ram_control[18]),.TB3S(GND),.C3Z(NET_356),.Q3Z(m1_ram_control[21]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_J16_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64_CAND2_TLSBR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T0I0(NET_627),.T0I1(NET_624),.T0I2(NET_626),.T0I3(NET_625),.TB0S(GND),.Q0Z(lint_RDATA_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J16_1 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64_CAND2_TLSBR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T1I0(NET_349),.T1I1(NET_351),.T1I2(NET_352),.T1I3(NET_350),.TB1S(GND),.Q1Z(lint_RDATA_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_J16_2 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0000000100000000),.B2I0(lint_ADDR_int[8]),.B2I1(lint_ADDR_int[7]),.B2I2(apb_fsm[0]),.B2I3(lint_ADDR_int[2]),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T2I0(GND),.T2I1(NET_336),.T2I2(NET_337),.T2I3(NET_338),.TB2S(GND),.B2Z(NET_10),.C2Z(NET_333),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J16_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF),.T3I0(NET_354),.T3I1(GND),.T3I2(NET_356),.T3I3(NET_355),.TB3S(GND),.C3Z(NET_352),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_J17_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_6),.B0I1(NET_5),.B0I2(fpgaio_out_dup_0[33]),.B0I3(tcdm_rdata_p2_int[1]),.CD0S(VCC),.Q0DI(lint_WDATA_int[17]),.Q0EN(nx19726z1_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T0I0(NET_6),.T0I1(NET_5),.T0I2(fpgaio_out_dup_0[41]),.T0I3(tcdm_rdata_p2_int[9]),.TB0S(GND),.B0Z(NET_2),.C0Z(NET_154),.Q0Z(m0_ram_control[17]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J17_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx19726z1_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p2_int[3]),.T1I1(NET_5),.T1I2(fpgaio_out_dup_0[35]),.T1I3(NET_6),.TB1S(GND),.C1Z(NET_688),.Q1Z(m0_ram_control[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_J17_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_94),.B2I1(m1_m0_dataout_int[17]),.B2I2(NET_103),.B2I3(m0_ram_control[17]),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p2_int[14]),.T2I1(NET_5),.T2I2(NET_6),.T2I3(fpgaio_out_dup_0[46]),.TB2S(GND),.B2Z(NET_337),.C2Z(NET_255),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J18_0 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_5),.B0I1(fpgaio_out_dup_0[47]),.B0I2(NET_6),.B0I3(tcdm_rdata_p2_int[15]),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.T0I0(NET_554),.T0I1(NET_555),.T0I2(NET_556),.T0I3(GND),.TB0S(GND),.B0Z(NET_294),.C0Z(NET_552),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J18_1 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.T1I0(GND),.T1I1(NET_409),.T1I2(NET_411),.T1I3(NET_410),.TB1S(GND),.C1Z(NET_407),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_J18_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.T2I0(NET_551),.T2I1(NET_549),.T2I2(NET_550),.T2I3(NET_552),.TB2S(GND),.Q2Z(lint_RDATA_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_J18_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.T3I0(NET_422),.T3I1(NET_423),.T3I2(NET_425),.T3I3(NET_424),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_J19_0 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_18_CAND5_BLSTR_10_tpGCLKBUF),.B0I1(m0_ram_control[27]),.B0I2(m1_m0_dataout_int[27]),.B0I3(NET_61),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx19726z1_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[11]),.T0I1(lint_ADDR_int[7]),.T0I2(NET_11),.T0I3(GND),.TB0S(GND),.B0Z(NET_546),.C0Z(NET_148),.Q0Z(m0_ram_control[27]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx19726z1_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q1Z(m0_ram_control[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J19_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T2I0(NET_31),.T2I1(GND),.T2I2(GND),.T2I3(NET_8),.TB2S(GND),.C2Z(NET_32),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J19_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_103),.T3I1(m1_m0_dataout_int[19]),.T3I2(m0_ram_control[19]),.T3I3(NET_94),.C3Z(NET_374),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J20_0 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_103),.B0I1(NET_94),.B0I2(m0_ram_control[21]),.B0I3(m1_m0_dataout_int[21]),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx19726z1_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[6]),.T0I1(NET_11),.T0I2(NET_10),.T0I3(lint_ADDR_int[5]),.TB0S(GND),.B0Z(NET_410),.C0Z(NET_17),.Q0Z(m0_ram_control[16]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_103),.B2I1(NET_94),.B2I2(m0_ram_control[18]),.B2I3(m1_m0_dataout_int[18]),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx19726z1_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B2Z(NET_355),.Q2Z(m0_ram_control[21]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J20_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx19726z1_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_61),.T3I1(NET_18_CAND5_BLSTR_10_tpGCLKBUF),.T3I2(m1_m0_dataout_int[16]),.T3I3(m0_ram_control[16]),.C3Z(NET_327),.Q3Z(m0_ram_control[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[17]),.Q0EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[49]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J21_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[8]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T1I0(m0_m0_dataout_int[20]),.T1I1(fpgaio_out_dup_0[52]),.T1I2(NET_59),.T1I3(NET_5),.C1Z(NET_392),.Q1Z(m1_m1_control[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J21_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_5),.B2I1(m0_m0_dataout_int[16]),.B2I2(fpgaio_out_dup_0[48]),.B2I3(NET_59),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T2I0(NET_29),.T2I1(NET_28_CAND4_BLSTR_10_tpGCLKBUF),.T2I2(m1_m1_control[8]),.T2I3(fpgaio_oe_dup_0[40]),.TB2S(GND),.B2Z(NET_317),.C2Z(NET_280),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx19726z1_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_rmode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J22_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T0I0(m1_ram_control[9]),.T0I1(NET_17_CAND3_BLSTR_10_tpGCLKBUF),.T0I2(m1_m0_dataout_int[9]),.T0I3(NET_18_CAND5_BLSTR_10_tpGCLKBUF),.TB0S(GND),.C0Z(NET_153),.Q0Z(fpgaio_out_dup_0[37]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_28_CAND4_BLSTR_10_tpGCLKBUF),.B2I1(NET_29),.B2I2(m1_m1_control[1]),.B2I3(fpgaio_oe_dup_0[33]),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B2Z(NET_25),.Q2Z(m1_ram_control[9]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J22_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_28_CAND4_BLSTR_10_tpGCLKBUF),.T3I1(NET_29),.T3I2(fpgaio_oe_dup_0[46]),.T3I3(m1_m1_osel_dup_0),.C3Z(NET_260),.Q3Z(m1_m1_control[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q0Z(m1_ram_control[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J23_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_17_CAND3_BLSTR_10_tpGCLKBUF),.T1I1(NET_18_CAND5_BLSTR_10_tpGCLKBUF),.T1I2(m1_m0_dataout_int[14]),.T1I3(m1_ram_control[14]),.TB1S(GND),.C1Z(NET_254),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_J23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_17_CAND3_BLSTR_10_tpGCLKBUF),.B2I1(NET_18_CAND5_BLSTR_10_tpGCLKBUF),.B2I2(m1_ram_control[15]),.B2I3(m1_m0_dataout_int[15]),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B2Z(NET_293),.Q2Z(m1_ram_control[15]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[58]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[50]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J29_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[9]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_32_CAND5_BLSBR_10_tpGCLKBUF),.T1I1(NET_33),.T1I2(m1_m1_dataout_int[9]),.T1I3(m1_m0_control[9]),.C1Z(NET_160),.Q1Z(m1_m0_control[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.Q3Z(m1_m0_outsel_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J30_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T0I0(m1_m1_dataout_int[14]),.T0I1(m1_m0_osel_dup_0),.T0I2(NET_33),.T0I3(NET_32_CAND5_BLSBR_10_tpGCLKBUF),.TB0S(GND),.C0Z(NET_261),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J30_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_dataout_int[4]),.T1I1(NET_33),.T1I2(m1_m0_outsel_dup_0[4]),.T1I3(NET_32_CAND5_BLSBR_10_tpGCLKBUF),.C1Z(NET_675),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J30_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T2I0(m1_m1_dataout_int[1]),.T2I1(NET_32_CAND5_BLSBR_10_tpGCLKBUF),.T2I2(m1_m0_outsel_dup_0[1]),.T2I3(NET_33),.TB2S(GND),.C2Z(NET_26),.Q2Z(m1_m0_outsel_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_J30_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_32_CAND5_BLSBR_10_tpGCLKBUF),.T3I1(m1_m1_dataout_int[3]),.T3I2(NET_33),.T3I3(m1_m0_outsel_dup_0[3]),.C3Z(NET_694),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J31_0 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1011101110110001),.B0I0(apb_fsm[0]),.B0I1(lint_ADDR_int[11]),.B0I2(lint_ADDR_int[13]),.B0I3(lint_ADDR_int[12]),.T0I0(apb_fsm[0]),.T0I1(lint_ADDR_int[11]),.T0I2(lint_ADDR_int[13]),.T0I3(lint_ADDR_int[12]),.TB0S(m1_oper0_rdata_int[20]),.C0Z(NET_745),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_J31_1 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1110000011101111),.B1I0(lint_ADDR_int[13]),.B1I1(lint_ADDR_int[12]),.B1I2(apb_fsm[0]),.B1I3(lint_ADDR_int[11]),.T1I0(apb_fsm[0]),.T1I1(lint_ADDR_int[11]),.T1I2(lint_ADDR_int[13]),.T1I3(lint_ADDR_int[12]),.TB1S(m1_oper0_rdata_int[16]),.C1Z(NET_743),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_J31_2 (.tFragBitInfo(16'b1011101110111011),.bFragBitInfo(16'b1011101110110001),.B2I0(apb_fsm[0]),.B2I1(lint_ADDR_int[11]),.B2I2(lint_ADDR_int[13]),.B2I3(lint_ADDR_int[12]),.T2I0(apb_fsm[0]),.T2I1(lint_ADDR_int[11]),.T2I2(lint_ADDR_int[13]),.T2I3(lint_ADDR_int[12]),.TB2S(m1_oper0_rdata_int[31]),.C2Z(NET_753),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_J31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K3_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_59),.B0I1(fpgaio_oe_dup_0[11]),.B0I2(m0_m0_dataout_int[11]),.B0I3(NET_58),.T0I0(NET_59),.T0I1(NET_58),.T0I2(fpgaio_oe_dup_0[5]),.T0I3(m0_m0_dataout_int[5]),.TB0S(GND),.B0Z(NET_209),.C0Z(NET_663),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K3_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B2I0(m0_m0_dataout_int[10]),.B2I1(fpgaio_oe_dup_0[10]),.B2I2(NET_59),.B2I3(NET_58),.T2I0(fpgaio_oe_dup_0[8]),.T2I1(m0_m0_dataout_int[8]),.T2I2(NET_59),.T2I3(NET_58),.TB2S(GND),.B2Z(NET_190),.C2Z(NET_289),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_K3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(NET_46_CAND1_TLSTR_11_tpGCLKBUF),.B3I1(NET_45),.B3I2(m0_oper1_rdata_int[8]),.B3I3(m1_oper0_rdata_int[8]),.T3I0(m0_oper1_rdata_int[8]),.T3I1(m1_oper0_rdata_int[8]),.T3I2(NET_46_CAND1_TLSTR_11_tpGCLKBUF),.T3I3(NET_45),.TB3S(NET_286),.C3Z(NET_284),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K4_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_58),.B0I1(NET_59),.B0I2(fpgaio_oe_dup_0[13]),.B0I3(m0_m0_dataout_int[13]),.T0I0(NET_59),.T0I1(fpgaio_oe_dup_0[4]),.T0I2(m0_m0_dataout_int[4]),.T0I3(NET_58),.TB0S(GND),.B0Z(NET_249),.C0Z(NET_683),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B1I0(m0_oper1_rdata_int[14]),.B1I1(m1_oper0_rdata_int[14]),.B1I2(NET_45),.B1I3(NET_46_CAND1_TLSTR_11_tpGCLKBUF),.T1I0(NET_45),.T1I1(NET_46_CAND1_TLSTR_11_tpGCLKBUF),.T1I2(m0_oper1_rdata_int[14]),.T1I3(m1_oper0_rdata_int[14]),.TB1S(NET_266),.C1Z(NET_264),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_K4_2 (.tFragBitInfo(16'b1010111110101111),.bFragBitInfo(16'b1010111110001101),.B2I0(apb_fsm[0]),.B2I1(lint_ADDR_int_13__CAND4_TLSTR_11_tpGCLKBUF),.B2I2(lint_ADDR_int[11]),.B2I3(lint_ADDR_int_14__CAND5_TLSTR_11_tpGCLKBUF),.T2I0(apb_fsm[0]),.T2I1(lint_ADDR_int_13__CAND4_TLSTR_11_tpGCLKBUF),.T2I2(lint_ADDR_int[11]),.T2I3(lint_ADDR_int_14__CAND5_TLSTR_11_tpGCLKBUF),.TB2S(m0_oper0_rdata_int[14]),.C2Z(NET_266),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_K4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(NET_46_CAND1_TLSTR_11_tpGCLKBUF),.B3I1(NET_45),.B3I2(m0_oper1_rdata_int[15]),.B3I3(m1_oper0_rdata_int[15]),.T3I0(m0_oper1_rdata_int[15]),.T3I1(m1_oper0_rdata_int[15]),.T3I2(NET_46_CAND1_TLSTR_11_tpGCLKBUF),.T3I3(NET_45),.TB3S(NET_305),.C3Z(NET_303),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(m0_oper1_rdata_int[3]),.B0I1(m1_oper0_rdata_int[3]),.B0I2(NET_46_CAND1_TLSTR_11_tpGCLKBUF),.B0I3(NET_45),.T0I0(m0_oper1_rdata_int[3]),.T0I1(m1_oper0_rdata_int[3]),.T0I2(NET_46_CAND1_TLSTR_11_tpGCLKBUF),.T0I3(NET_45),.TB0S(NET_699),.C0Z(NET_697),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_45),.B2I1(m1_oper0_rdata_int[4]),.B2I2(NET_46_CAND1_TLSTR_11_tpGCLKBUF),.B2I3(m0_oper1_rdata_int[4]),.T2I0(NET_45),.T2I1(m1_oper0_rdata_int[4]),.T2I2(NET_46_CAND1_TLSTR_11_tpGCLKBUF),.T2I3(m0_oper1_rdata_int[4]),.TB2S(NET_680),.C2Z(NET_678),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_K5_3 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int_14__CAND5_TLSTR_11_tpGCLKBUF),.T3I1(lint_ADDR_int[12]),.T3I2(apb_fsm[0]),.T3I3(GND),.TB3S(GND),.C3Z(NET_46),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m0_coef_rmode_dup_0[0]),.B0I1(NET_61),.B0I2(fpgaio_out_dup_0[8]),.B0I3(NET_60),.B0Z(NET_290),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K7_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_287),.B2I1(NET_290),.B2I2(NET_289),.B2I3(NET_288),.T2I0(NET_682),.T2I1(NET_684),.T2I2(NET_683),.T2I3(NET_681),.TB2S(GND),.B2Z(NET_291),.C2Z(NET_685),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_K7_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(fpgaio_out_dup_0[14]),.T3I1(NET_61),.T3I2(NET_60),.T3I3(m0_coef_wdsel_dup_0),.TB3S(GND),.C3Z(NET_270),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K8_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_61),.T1I1(fpgaio_out_dup_0[11]),.T1I2(m0_coef_wmode_dup_0[1]),.T1I3(NET_60),.TB1S(GND),.C1Z(NET_210),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_K8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K8_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_191),.T3I1(NET_189),.T3I2(NET_190),.T3I3(NET_188),.TB3S(GND),.C3Z(NET_192),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K9_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.T0I0(m0_m1_outsel_dup_0[2]),.T0I1(NET_111),.T0I2(fpgaio_in_int[2]),.T0I3(NET_112),.TB0S(GND),.C0Z(NET_717),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K9_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_210),.T1I1(NET_207),.T1I2(NET_209),.T1I3(NET_208),.TB1S(GND),.C1Z(NET_211),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_K9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_111),.B2I1(m0_m1_outsel_dup_0[0]),.B2I2(fpgaio_in_int[0]),.B2I3(NET_112),.B2Z(NET_107),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K9_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(fpgaio_in_int[6]),.T3I1(NET_111),.T3I2(m0_m1_tc_dup_0),.T3I3(NET_112),.TB3S(GND),.C3Z(NET_636),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K10_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_in_int[7]),.B0I1(NET_112),.B0I2(NET_111),.B0I3(m0_m1_control[7]),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(NET_111),.T0I1(NET_112),.T0I2(m0_m1_mode_dup_0[0]),.T0I3(fpgaio_in_int[12]),.TB0S(GND),.B0Z(NET_470),.C0Z(NET_224),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K10_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_13),.T1I1(tcdm_result_p0[4]),.T1I2(NET_12),.T1I3(fpgaio_out_dup_0[68]),.C1Z(NET_670),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K10_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_13),.T2I1(fpgaio_out_dup_0[69]),.T2I2(NET_12),.T2I3(tcdm_result_p0[5]),.TB2S(GND),.C2Z(NET_650),.Q2Z(m0_m0_outsel_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_K10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_mode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_13),.B0I1(fpgaio_out_dup_0[74]),.B0I2(tcdm_result_p0[10]),.B0I3(NET_12),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.B0Z(NET_177),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K11_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T1I0(NET_13),.T1I1(NET_12),.T1I2(tcdm_result_p0[11]),.T1I3(fpgaio_out_dup_0[75]),.TB1S(GND),.C1Z(NET_196),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_K11_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_13),.B2I1(NET_12),.B2I2(tcdm_result_p0[13]),.B2I3(fpgaio_out_dup_0[77]),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T2I0(NET_13),.T2I1(fpgaio_out_dup_0[72]),.T2I2(NET_12),.T2I3(tcdm_result_p0[8]),.TB2S(GND),.B2Z(NET_236),.C2Z(NET_276),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K11_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_740),.B3I1(NET_282),.B3I2(NET_285),.B3I3(NET_277),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64_CAND2_TLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T3I0(NET_285),.T3I1(NET_277),.T3I2(NET_740),.T3I3(NET_282),.TB3S(NET_291),.Q3Z(lint_RDATA_dup_0[8]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_K12_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(GND),.B0I1(RESET_int[0]),.B0I2(GND),.B0I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T0I0(NET_193),.T0I1(NET_195),.T0I2(NET_194),.T0I3(NET_196),.TB0S(GND),.B0Z(not_RESET_0),.C0Z(NET_197),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K12_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T1I0(NET_275),.T1I1(NET_276),.T1I2(NET_274),.T1I3(NET_273),.TB1S(GND),.C1Z(NET_277),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_K12_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_205),.B2I1(NET_734),.B2I2(NET_202),.B2I3(NET_197),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64_CAND2_TLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T2I0(NET_205),.T2I1(NET_734),.T2I2(NET_202),.T2I3(NET_197),.TB2S(NET_211),.Q2Z(lint_RDATA_dup_0[11]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_K12_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T3I0(NET_235),.T3I1(NET_233),.T3I2(NET_236),.T3I3(NET_234),.TB3S(GND),.C3Z(NET_237),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_K13_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_676),.B0I1(NET_759),.B0I2(NET_671),.B0I3(NET_679),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z64_CAND2_TLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T0I0(NET_676),.T0I1(NET_759),.T0I2(NET_671),.T0I3(NET_679),.TB0S(NET_685),.Q0Z(lint_RDATA_dup_0[4]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K13_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T1I0(NET_668),.T1I1(NET_669),.T1I2(NET_667),.T1I3(NET_670),.TB1S(GND),.C1Z(NET_671),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_K13_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T2I0(NET_201),.T2I1(NET_198),.T2I2(NET_200),.T2I3(NET_199),.TB2S(GND),.C2Z(NET_202),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K13_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_304),.B3I1(NET_301),.B3I2(NET_742),.B3I3(NET_296),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64_CAND2_TLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T3I0(NET_742),.T3I1(NET_296),.T3I2(NET_304),.T3I3(NET_301),.TB3S(NET_310),.Q3Z(lint_RDATA_dup_0[15]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_K14_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_175),.B0I1(NET_176),.B0I2(NET_177),.B0I3(NET_174),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T0I0(NET_179),.T0I1(NET_181),.T0I2(NET_182),.T0I3(NET_180),.TB0S(GND),.B0Z(NET_178),.C0Z(NET_183),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_300),.B2I1(NET_299),.B2I2(NET_297),.B2I3(NET_298),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.B2Z(NET_301),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K14_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_178),.B3I1(NET_183),.B3I2(NET_186),.B3I3(NET_732),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64_CAND2_TLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T3I0(NET_186),.T3I1(NET_732),.T3I2(NET_178),.T3I3(NET_183),.TB3S(NET_192),.Q3Z(lint_RDATA_dup_0[10]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_K15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_104),.B0I1(NET_107),.B0I2(NET_106),.B0I3(NET_105),.B0Z(NET_79),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K15_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_468),.T1I1(NET_469),.T1I2(NET_467),.T1I3(NET_470),.TB1S(GND),.C1Z(NET_459),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_K15_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_279),.B2I1(NET_278),.B2I2(NET_280),.B2I3(NET_281),.T2I0(NET_222),.T2I1(NET_221),.T2I2(NET_223),.T2I3(NET_224),.TB2S(GND),.B2Z(NET_282),.C2Z(NET_213),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_K15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K16_0 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T0I0(GND),.T0I1(NET_373),.T0I2(NET_375),.T0I3(NET_374),.TB0S(GND),.C0Z(NET_371),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K16_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T1I0(NET_633),.T1I1(NET_635),.T1I2(NET_634),.T1I3(NET_636),.TB1S(GND),.C1Z(NET_625),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_K16_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64_CAND2_TLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T2I0(NET_332),.T2I1(NET_331),.T2I2(NET_330),.T2I3(NET_333),.TB2S(GND),.Q2Z(lint_RDATA_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_K16_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64_CAND2_TLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF),.T3I0(NET_370),.T3I1(NET_369),.T3I2(NET_368),.T3I3(NET_371),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_K17_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B0I0(tcdm_rdata_p2_int[11]),.B0I1(fpgaio_out_dup_0[43]),.B0I2(NET_5),.B0I3(NET_6),.T0I0(fpgaio_out_dup_0[42]),.T0I1(NET_6),.T0I2(tcdm_rdata_p2_int[10]),.T0I3(NET_5),.TB0S(GND),.B0Z(NET_195),.C0Z(NET_176),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K17_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_717),.T2I1(NET_716),.T2I2(NET_715),.T2I3(NET_714),.TB2S(GND),.C2Z(NET_706),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_K17_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(tcdm_rdata_p2_int[5]),.T3I1(fpgaio_out_dup_0[37]),.T3I2(NET_6),.T3I3(NET_5),.TB3S(GND),.C3Z(NET_649),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K18_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.T0I0(tcdm_rdata_p2_int[4]),.T0I1(NET_6),.T0I2(NET_5),.T0I3(fpgaio_out_dup_0[36]),.TB0S(GND),.C0Z(NET_669),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K18_1 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.T1I0(NET_407),.T1I1(NET_405),.T1I2(NET_406),.T1I3(NET_404),.TB1S(GND),.Q1Z(lint_RDATA_dup_0[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_K18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(fpgaio_out_dup_0[40]),.B2I1(NET_6),.B2I2(NET_5),.B2I3(tcdm_rdata_p2_int[8]),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.B2Z(NET_275),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K18_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.T3I0(NET_6),.T3I1(NET_5),.T3I2(fpgaio_out_dup_0[45]),.T3I3(tcdm_rdata_p2_int[13]),.TB3S(GND),.C3Z(NET_235),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_K19_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000010000000),.B0I0(NET_71),.B0I1(NET_73),.B0I2(NET_72),.B0I3(GND),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx19726z1_CAND2_BLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T0I0(NET_18_CAND5_BLSTR_11_tpGCLKBUF),.T0I1(NET_61),.T0I2(m0_ram_control[30]),.T0I3(m1_m0_dataout_int[30]),.TB0S(GND),.B0Z(NET_69),.C0Z(NET_599),.Q0Z(m0_ram_control[20]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K19_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_148),.T1I1(NET_602),.T1I2(NET_70),.T1I3(NET_69),.TB1S(GND),.C1Z(nx4939z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_K19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B2I0(NET_148),.B2I1(GND),.B2I2(GND),.B2I3(NET_69),.CD2S(VCC),.Q2DI(lint_WDATA_int[30]),.Q2EN(nx19726z1_CAND2_BLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.B2Z(NET_146),.Q2Z(m0_ram_control[30]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K19_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(m0_ram_control[20]),.T3I1(NET_61),.T3I2(m1_m0_dataout_int[20]),.T3I3(NET_18_CAND5_BLSTR_11_tpGCLKBUF),.C3Z(NET_401),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_K20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000010),.B0I0(apb_fsm[0]),.B0I1(apb_fsm[1]),.B0I2(GND),.B0I3(GND),.B0Z(NET_65),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K20_1 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[15]),.T1I1(lint_ADDR_int[12]),.T1I2(lint_ADDR_int[14]),.T1I3(NET_73),.C1Z(NET_149),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000100000000),.B2I0(lint_ADDR_int[15]),.B2I1(lint_ADDR_int[10]),.B2I2(lint_ADDR_int[8]),.B2I3(NET_74),.B2Z(NET_72),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K20_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int[13]),.T3I1(lint_ADDR_int[12]),.T3I2(lint_ADDR_int[14]),.T3I3(GND),.TB3S(GND),.C3Z(NET_74),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_K21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q0Z(m1_ram_control[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[43]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K21_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T2I0(m1_ram_control[11]),.T2I1(m1_m0_dataout_int[11]),.T2I2(NET_18_CAND5_BLSTR_11_tpGCLKBUF),.T2I3(NET_17_CAND3_BLSTR_11_tpGCLKBUF),.TB2S(GND),.C2Z(NET_194),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K21_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_dataout_int[8]),.T3I1(NET_18_CAND5_BLSTR_11_tpGCLKBUF),.T3I2(m1_ram_control[8]),.T3I3(NET_17_CAND3_BLSTR_11_tpGCLKBUF),.C3Z(NET_274),.Q3Z(m1_ram_control[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_K22_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T0I0(NET_18_CAND5_BLSTR_11_tpGCLKBUF),.T0I1(m1_m0_dataout_int[10]),.T0I2(NET_17_CAND3_BLSTR_11_tpGCLKBUF),.T0I3(m1_ram_control[10]),.TB0S(GND),.C0Z(NET_175),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K22_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_oe_dup_0[47]),.T1I1(NET_28_CAND4_BLSTR_11_tpGCLKBUF),.T1I2(m1_m1_csel_dup_0),.T1I3(NET_29),.TB1S(GND),.C1Z(NET_299),.Q1Z(m1_ram_control[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_K22_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_m1_mode_dup_0[1]),.B2I1(NET_28_CAND4_BLSTR_11_tpGCLKBUF),.B2I2(fpgaio_oe_dup_0[45]),.B2I3(NET_29),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_317),.T2I1(NET_320),.T2I2(NET_319),.T2I3(NET_318),.TB2S(GND),.B2Z(NET_240),.C2Z(NET_314),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K23_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T0I0(m1_m0_dataout_int[13]),.T0I1(NET_18_CAND5_BLSTR_11_tpGCLKBUF),.T0I2(m1_ram_control[13]),.T0I3(NET_17_CAND3_BLSTR_11_tpGCLKBUF),.TB0S(GND),.C0Z(NET_234),.Q0Z(fpgaio_out_dup_0[55]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K23_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_17_CAND3_BLSTR_11_tpGCLKBUF),.T1I1(NET_18_CAND5_BLSTR_11_tpGCLKBUF),.T1I2(m1_ram_control[1]),.T1I3(m1_m0_dataout_int[1]),.TB1S(GND),.C1Z(NET_1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_K23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q2Z(m1_ram_control[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q3Z(m1_ram_control[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q3Z(m1_m0_tc_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K30_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B0I0(m1_m0_csel_dup_0),.B0I1(NET_33),.B0I2(m1_m1_dataout_int[15]),.B0I3(NET_32_CAND5_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(NET_32_CAND5_BLSBR_11_tpGCLKBUF),.T0I1(NET_33),.T0I2(m1_m0_control[11]),.T0I3(m1_m1_dataout_int[11]),.TB0S(GND),.B0Z(NET_300),.C0Z(NET_201),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_csel_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K30_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(NET_32_CAND5_BLSBR_11_tpGCLKBUF),.T3I1(NET_33),.T3I2(m1_m0_rnd_dup_0),.T3I3(m1_m1_dataout_int[16]),.C3Z(NET_318),.Q3Z(m1_m0_control[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_K31_0 (.tFragBitInfo(16'b1111111100110011),.bFragBitInfo(16'b1111101000110011),.B0I0(lint_ADDR_int[12]),.B0I1(lint_ADDR_int[11]),.B0I2(lint_ADDR_int[13]),.B0I3(apb_fsm[0]),.T0I0(lint_ADDR_int[12]),.T0I1(lint_ADDR_int[11]),.T0I2(lint_ADDR_int[13]),.T0I3(apb_fsm[0]),.TB0S(m1_oper0_rdata_int[30]),.C0Z(NET_751),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K32_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_43_CAND3_BLSBR_11_tpGCLKBUF),.B0I1(m1_coef_rdata_int[24]),.B0I2(m1_oper0_rdata_int[24]),.B0I3(NET_45),.T0I0(m1_coef_rdata_int[28]),.T0I1(m1_oper0_rdata_int[28]),.T0I2(NET_43_CAND3_BLSBR_11_tpGCLKBUF),.T0I3(NET_45),.TB0S(GND),.B0Z(NET_494),.C0Z(NET_564),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_K32_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_43_CAND3_BLSBR_11_tpGCLKBUF),.T1I1(m1_oper0_rdata_int[26]),.T1I2(m1_coef_rdata_int[26]),.T1I3(NET_45),.C1Z(NET_529),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K32_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m1_coef_rdata_int[29]),.T3I1(NET_43_CAND3_BLSBR_11_tpGCLKBUF),.T3I2(m1_oper0_rdata_int[29]),.T3I3(NET_45),.TB3S(GND),.C3Z(NET_582),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_L1_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B0I0(m0_oper0_rdata_int[7]),.B0I1(NET_117),.B0I2(m0_oper1_rdata_int[7]),.B0I3(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.T0I0(m0_oper1_rdata_int[2]),.T0I1(m0_oper0_rdata_int[2]),.T0I2(NET_117),.T0I3(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.TB0S(GND),.B0Z(NET_472),.C0Z(NET_719),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_L1_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_oper0_rdata_int[6]),.T1I1(NET_117),.T1I2(m0_oper1_rdata_int[6]),.T1I3(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.C1Z(NET_638),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_L1_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.B2I1(NET_117),.B2I2(m0_oper0_rdata_int[12]),.B2I3(m0_oper1_rdata_int[12]),.T2I0(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.T2I1(NET_117),.T2I2(m0_oper0_rdata_int[0]),.T2I3(m0_oper1_rdata_int[0]),.TB2S(GND),.B2Z(NET_226),.C2Z(NET_114),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_L1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.B0I1(m0_oper1_rdata_int[13]),.B0I2(NET_45),.B0I3(m1_oper0_rdata_int[13]),.T0I0(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.T0I1(m0_oper1_rdata_int[13]),.T0I2(NET_45),.T0I3(m1_oper0_rdata_int[13]),.TB0S(NET_246),.C0Z(NET_244),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_L3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(NET_45),.B1I1(m1_oper0_rdata_int[9]),.B1I2(m0_oper1_rdata_int[9]),.B1I3(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.T1I0(m0_oper1_rdata_int[9]),.T1I1(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.T1I2(NET_45),.T1I3(m1_oper0_rdata_int[9]),.TB1S(NET_165),.C1Z(NET_163),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_L3_2 (.tFragBitInfo(16'b0100110000000000),.bFragBitInfo(16'b0111000000000000),.B2I0(m0_coef_rdata_int[8]),.B2I1(NET_41),.B2I2(NET_284),.B2I3(NET_283),.T2I0(NET_41),.T2I1(NET_162),.T2I2(m0_coef_rdata_int[9]),.T2I3(NET_163),.TB2S(GND),.B2Z(NET_285),.C2Z(NET_164),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_L3_3 (.tFragBitInfo(16'b0000100010001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_244),.T3I1(NET_243),.T3I2(NET_41),.T3I3(m0_coef_rdata_int[13]),.C3Z(NET_245),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.B0I1(m1_oper0_rdata_int[10]),.B0I2(NET_45),.B0I3(m0_oper1_rdata_int[10]),.T0I0(NET_46_CAND1_TLSTR_12_tpGCLKBUF),.T0I1(m1_oper0_rdata_int[10]),.T0I2(NET_45),.T0I3(m0_oper1_rdata_int[10]),.TB0S(NET_187),.C0Z(NET_185),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_L4_1 (.tFragBitInfo(16'b1010111110101111),.bFragBitInfo(16'b1111010111000101),.B1I0(lint_ADDR_int[11]),.B1I1(lint_ADDR_int_14__CAND5_TLSTR_12_tpGCLKBUF),.B1I2(apb_fsm[0]),.B1I3(lint_ADDR_int_13__CAND4_TLSTR_12_tpGCLKBUF),.T1I0(apb_fsm[0]),.T1I1(lint_ADDR_int_13__CAND4_TLSTR_12_tpGCLKBUF),.T1I2(lint_ADDR_int[11]),.T1I3(lint_ADDR_int_14__CAND5_TLSTR_12_tpGCLKBUF),.TB1S(m0_oper0_rdata_int[10]),.C1Z(NET_187),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_L4_2 (.tFragBitInfo(16'b0111000000000000),.bFragBitInfo(16'b0010000010100000),.B2I0(NET_185),.B2I1(m0_coef_rdata_int[10]),.B2I2(NET_184),.B2I3(NET_41),.T2I0(NET_41),.T2I1(m0_coef_rdata_int[14]),.T2I2(NET_264),.T2I3(NET_263),.TB2S(GND),.B2Z(NET_186),.C2Z(NET_265),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_L4_3 (.tFragBitInfo(16'b0100110000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m0_coef_rdata_int[15]),.T3I1(NET_302),.T3I2(NET_41),.T3I3(NET_303),.C3Z(NET_304),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L7_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[9]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND3_TLSTR_12_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_out_dup_0[4]),.T0I1(m0_oper1_rmode_dup_0[0]),.T0I2(NET_60),.T0I3(NET_61),.TB0S(GND),.C0Z(NET_684),.Q0Z(tcdm_result_p0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L7_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND3_TLSTR_12_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[13]),.T1I1(NET_61),.T1I2(NET_60),.T1I3(m0_oper1_wdsel_dup_0),.TB1S(GND),.C1Z(NET_250),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L7_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_60),.B2I1(m0_oper1_rmode_dup_0[1]),.B2I2(fpgaio_out_dup_0[5]),.B2I3(NET_61),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND3_TLSTR_12_tpGCLKBUF),.QST(GND),.T2I0(NET_661),.T2I1(NET_663),.T2I2(NET_664),.T2I3(NET_662),.TB2S(GND),.B2Z(NET_664),.C2Z(NET_665),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_L7_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[8]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND3_TLSTR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_248),.T3I1(NET_247),.T3I2(NET_249),.T3I3(NET_250),.TB3S(GND),.C3Z(NET_251),.Q3Z(tcdm_result_p0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L8_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B0I0(tcdm_result_p0[6]),.B0I1(NET_89),.B0I2(m0_m0_dataout_int[6]),.B0I3(NET_95),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[7]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND3_TLSTR_12_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p0[6]),.T0I1(NET_89),.T0I2(m0_m0_dataout_int[6]),.T0I3(NET_95),.TB0S(NET_15),.C0Z(NET_637),.Q0Z(tcdm_result_p0[7]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L8_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(tcdm_result_p0[2]),.B1I1(NET_95),.B1I2(NET_89),.B1I3(m0_m0_dataout_int[2]),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND3_TLSTR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_89),.T1I1(m0_m0_dataout_int[2]),.T1I2(tcdm_result_p0[2]),.T1I3(NET_95),.TB1S(NET_15),.C1Z(NET_718),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L8_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[6]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND3_TLSTR_12_tpGCLKBUF),.QST(GND),.T2I0(m0_coef_wmode_dup_0[0]),.T2I1(NET_60),.T2I2(fpgaio_out_dup_0[10]),.T2I3(NET_61),.TB2S(GND),.C2Z(NET_191),.Q2Z(tcdm_result_p0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_L8_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B3I0(m0_m0_dataout_int[7]),.B3I1(NET_95),.B3I2(tcdm_result_p0[7]),.B3I3(NET_89),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[2]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND3_TLSTR_12_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p0[7]),.T3I1(NET_89),.T3I2(m0_m0_dataout_int[7]),.T3I3(NET_95),.TB3S(NET_15),.C3Z(NET_471),.Q3Z(tcdm_result_p0[2]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L9_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B0I0(tcdm_result_p0[0]),.B0I1(NET_89),.B0I2(NET_95),.B0I3(m0_m0_dataout_int[0]),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[12]),.Q0EN(tcdm_valid_p0_int_CAND1_TLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p0[0]),.T0I1(NET_89),.T0I2(NET_95),.T0I3(m0_m0_dataout_int[0]),.TB0S(NET_15_CAND5_TLSBR_12_tpGCLKBUF),.C0Z(NET_113),.Q0Z(tcdm_result_p0[12]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L9_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(m1_coef_rdata_int[12]),.T1I1(NET_43),.T1I2(m0_coef_rdata_int[12]),.T1I3(NET_41),.TB1S(GND),.C1Z(NET_227),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_228),.B2I1(NET_225),.B2I2(NET_226),.B2I3(NET_227),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[0]),.Q2EN(tcdm_valid_p0_int_CAND1_TLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.B2Z(NET_222),.Q2Z(tcdm_result_p0[0]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L9_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B3I0(NET_95),.B3I1(m0_m0_dataout_int[12]),.B3I2(tcdm_result_p0[12]),.B3I3(NET_89),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[3]),.Q3EN(tcdm_valid_p0_int_CAND1_TLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p0[12]),.T3I1(NET_89),.T3I2(NET_95),.T3I3(m0_m0_dataout_int[12]),.TB3S(NET_15_CAND5_TLSBR_12_tpGCLKBUF),.C3Z(NET_225),.Q3Z(tcdm_result_p0[3]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L10_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(NET_639),.T0I1(NET_638),.T0I2(NET_640),.T0I3(NET_637),.TB0S(GND),.C0Z(NET_634),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L10_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_721),.T1I1(NET_719),.T1I2(NET_718),.T1I3(NET_720),.TB1S(GND),.C1Z(NET_715),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_116),.B2I1(NET_114),.B2I2(NET_115),.B2I3(NET_113),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.B2Z(NET_105),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L10_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_472),.T3I1(NET_471),.T3I2(NET_474),.T3I3(NET_473),.TB3S(GND),.C3Z(NET_468),.Q3Z(m0_m1_control[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(lint_ADDR_int[11]),.B0I1(lint_ADDR_int[2]),.B0I2(lint_ADDR_int[7]),.B0I3(apb_fsm[0]),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[11]),.T0I1(lint_ADDR_int[2]),.T0I2(lint_ADDR_int[7]),.T0I3(apb_fsm[0]),.TB0S(lint_ADDR_int[8]),.C0Z(NET_95),.Q0Z(m0_m0_outsel_dup_0[5]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L12_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.T0I0(NET_655),.T0I1(NET_652),.T0I2(NET_653),.T0I3(NET_654),.TB0S(GND),.C0Z(NET_656),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L12_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B1I0(NET_651),.B1I1(NET_656),.B1I2(NET_757),.B1I3(NET_659),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64_CAND2_TLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.T1I0(NET_757),.T1I1(NET_659),.T1I2(NET_651),.T1I3(NET_656),.TB1S(NET_665),.Q1Z(lint_RDATA_dup_0[5]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_L12_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_237),.B2I1(NET_242),.B2I2(NET_736),.B2I3(NET_245),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64_CAND2_TLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.T2I0(NET_237),.T2I1(NET_242),.T2I2(NET_736),.T2I3(NET_245),.TB2S(NET_251),.Q2Z(lint_RDATA_dup_0[13]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_L12_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.T3I0(NET_650),.T3I1(NET_648),.T3I2(NET_647),.T3I3(NET_649),.C3Z(NET_651),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L14_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.T0I0(NET_240),.T0I1(NET_238),.T0I2(NET_241),.T0I3(NET_239),.TB0S(GND),.C0Z(NET_242),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_L14_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_oper0_rdata_int[21]),.T1I1(NET_44),.T1I2(m1_oper1_rdata_int[21]),.T1I3(NET_117),.TB1S(GND),.C1Z(NET_420),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_L14_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000001000000),.B2I0(lint_ADDR_int[7]),.B2I1(NET_19),.B2I2(NET_15_CAND5_TLSBR_12_tpGCLKBUF),.B2I3(lint_ADDR_int[2]),.T2I0(m1_oper1_rdata_int[29]),.T2I1(NET_44),.T2I2(NET_117),.T2I3(m0_oper0_rdata_int[29]),.TB2S(GND),.B2Z(NET_59),.C2Z(NET_583),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_L14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100010001000),.B3I0(NET_419),.B3I1(NET_420),.B3I2(NET_124_CAND4_TLSBR_12_tpGCLKBUF),.B3I3(tcdm_rdata_p0_int[21]),.T3I0(NET_124_CAND4_TLSBR_12_tpGCLKBUF),.T3I1(tcdm_rdata_p0_int[21]),.T3I2(NET_419),.T3I3(NET_420),.TB3S(NET_421),.C3Z(NET_404),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_L15_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000001000000000),.B0I0(NET_95),.B0I1(GND),.B0I2(GND),.B0I3(NET_15_CAND5_TLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(m0_oper0_rdata_int[26]),.T0I1(NET_117),.T0I2(m1_oper1_rdata_int[26]),.T0I3(NET_44),.TB0S(GND),.B0Z(NET_334),.C0Z(NET_530),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L15_1 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_95),.T1I1(GND),.T1I2(GND),.T1I3(NET_7),.TB1S(GND),.C1Z(NET_94),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010101000000000),.B2I0(NET_530),.B2I1(NET_124_CAND4_TLSBR_12_tpGCLKBUF),.B2I2(tcdm_rdata_p0_int[26]),.B2I3(NET_529),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T2I0(NET_530),.T2I1(NET_124_CAND4_TLSBR_12_tpGCLKBUF),.T2I2(tcdm_rdata_p0_int[26]),.T2I3(NET_529),.TB2S(NET_531),.C2Z(NET_514),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_L15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010101000000000),.B3I0(NET_582),.B3I1(NET_124_CAND4_TLSBR_12_tpGCLKBUF),.B3I2(tcdm_rdata_p0_int[29]),.B3I3(NET_583),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p0_int[29]),.T3I1(NET_583),.T3I2(NET_582),.T3I3(NET_124_CAND4_TLSBR_12_tpGCLKBUF),.TB3S(NET_584),.C3Z(NET_567),.Q3Z(m0_m0_outsel_dup_0[2]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_334),.B0I1(tcdm_result_p2[17]),.B0I2(m0_m0_dataout_int[17]),.B0I3(NET_82),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(NET_334),.T0I1(tcdm_result_p2[17]),.T0I2(m0_m0_dataout_int[17]),.T0I3(NET_82),.TB0S(NET_335),.C0Z(NET_332),.Q0Z(m0_m0_control[7]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(tcdm_result_p2[19]),.B1I1(NET_82),.B1I2(NET_334),.B1I3(m0_m0_dataout_int[19]),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_334),.T1I1(m0_m0_dataout_int[19]),.T1I2(tcdm_result_p2[19]),.T1I3(NET_82),.TB1S(NET_372),.C1Z(NET_370),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_334),.B2I1(m0_m0_dataout_int[18]),.B2I2(tcdm_result_p2[18]),.B2I3(NET_82),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T2I0(NET_334),.T2I1(m0_m0_dataout_int[18]),.T2I2(tcdm_result_p2[18]),.T2I3(NET_82),.TB2S(NET_353),.C2Z(NET_351),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_L16_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[19]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p2_int[7]),.T3I1(NET_109),.T3I2(NET_108),.T3I3(m0_m0_control[7]),.C3Z(NET_469),.Q3Z(tcdm_result_p2[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L17_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p2_int[22]),.T0I1(NET_109),.T0I2(m0_m1_control[22]),.T0I3(NET_112),.TB0S(GND),.C0Z(NET_433),.Q0Z(m0_m1_control[29]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B1I0(tcdm_result_p2[22]),.B1I1(NET_334),.B1I2(NET_82),.B1I3(m0_m0_dataout_int[22]),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[22]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_82),.T1I1(m0_m0_dataout_int[22]),.T1I2(tcdm_result_p2[22]),.T1I3(NET_334),.TB1S(NET_426),.C1Z(NET_424),.Q1Z(tcdm_result_p2[22]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_L17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_82),.B2I1(tcdm_result_p2[29]),.B2I2(NET_334),.B2I3(m0_m0_dataout_int[29]),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[29]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T2I0(NET_82),.T2I1(tcdm_result_p2[29]),.T2I2(NET_334),.T2I3(m0_m0_dataout_int[29]),.TB2S(NET_571),.C2Z(NET_569),.Q2Z(tcdm_result_p2[29]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_L17_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T3I0(m0_m1_control[29]),.T3I1(NET_109),.T3I2(tcdm_rdata_p2_int[29]),.T3I3(NET_112),.TB3S(GND),.C3Z(NET_578),.Q3Z(m0_m1_control[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(tcdm_rdata_p2_int[26]),.B0I1(NET_109),.B0I2(NET_112),.B0I3(m0_m1_control[26]),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[24]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B0Z(NET_525),.Q0Z(tcdm_result_p2[24]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(NET_334),.B1I1(m0_m0_dataout_int[24]),.B1I2(tcdm_result_p2[24]),.B1I3(NET_82),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[21]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p2[24]),.T1I1(NET_82),.T1I2(NET_334),.T1I3(m0_m0_dataout_int[24]),.TB1S(NET_483),.C1Z(NET_481),.Q1Z(tcdm_result_p2[21]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_L18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m0_m1_control[21]),.B2I1(NET_109),.B2I2(NET_112),.B2I3(tcdm_rdata_p2_int[21]),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B2Z(NET_415),.Q2Z(m0_m1_control[21]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(NET_334),.B3I1(tcdm_result_p2[21]),.B3I2(m0_m0_dataout_int[21]),.B3I3(NET_82),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_dataout_int[21]),.T3I1(NET_82),.T3I2(NET_334),.T3I3(tcdm_result_p2[21]),.TB3S(NET_408),.C3Z(NET_406),.Q3Z(m0_m1_control[26]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L19_0 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[2]),.T0I1(NET_19),.T0I2(lint_ADDR_int[7]),.T0I3(NET_7),.TB0S(GND),.C0Z(NET_18),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L19_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx19726z1_CAND2_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[4]),.T1I1(NET_69),.T1I2(NET_70),.T1I3(GND),.TB1S(GND),.C1Z(NET_67),.Q1Z(m0_oper1_wdsel_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_L19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L19_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx19726z1_CAND2_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_18_CAND5_BLSTR_12_tpGCLKBUF),.T3I1(NET_61),.T3I2(m1_m0_dataout_int[31]),.T3I3(m0_ram_control[31]),.TB3S(GND),.C3Z(NET_617),.Q3Z(m0_ram_control[31]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx19726z1_CAND2_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wmode_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L20_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T1I0(m1_m0_dataout_int[3]),.T1I1(NET_17_CAND3_BLSTR_12_tpGCLKBUF),.T1I2(m1_ram_control[3]),.T1I3(NET_18_CAND5_BLSTR_12_tpGCLKBUF),.TB1S(GND),.C1Z(NET_687),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(m1_ram_control[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L20_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx19726z1_CAND2_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_18_CAND5_BLSTR_12_tpGCLKBUF),.T3I1(m1_m0_dataout_int[25]),.T3I2(NET_61),.T3I3(m0_ram_control[25]),.TB3S(GND),.C3Z(NET_511),.Q3Z(m0_ram_control[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_L22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_m1_osel_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx19726z1_CAND2_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_rmode_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx19726z1_CAND2_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_rmode_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_csel_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_control[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L23_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T1I0(m1_m0_dataout_int[4]),.T1I1(NET_17_CAND3_BLSTR_12_tpGCLKBUF),.T1I2(m1_ram_control[4]),.T1I3(NET_18_CAND5_BLSTR_12_tpGCLKBUF),.TB1S(GND),.C1Z(NET_668),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(m1_m0_dataout_int[5]),.B2I1(NET_17_CAND3_BLSTR_12_tpGCLKBUF),.B2I2(m1_ram_control[5]),.B2I3(NET_18_CAND5_BLSTR_12_tpGCLKBUF),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B2Z(NET_648),.Q2Z(m1_ram_control[5]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L23_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T3I0(m1_m1_dataout_int[8]),.T3I1(m1_m0_control[8]),.T3I2(NET_32),.T3I3(NET_33),.C3Z(NET_281),.Q3Z(m1_ram_control[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L27_3 (.tFragBitInfo(16'b0000000000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(apb_fsm[0]),.T3I1(lint_ADDR_int[13]),.T3I2(lint_ADDR_int[12]),.T3I3(GND),.C3Z(NET_45),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L30_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_33),.T3I1(m1_m0_outsel_dup_0[5]),.T3I2(m1_m1_dataout_int[5]),.T3I3(NET_32_CAND5_BLSBR_12_tpGCLKBUF),.TB3S(GND),.C3Z(NET_655),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_L31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L31_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m1_oper0_rdata_int[2]),.T1I1(m1_oper1_rdata_int[2]),.T1I2(NET_45),.T1I3(NET_44_CAND4_BLSBR_12_tpGCLKBUF),.TB1S(GND),.C1Z(NET_721),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_L31_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.T2I0(m1_oper0_rdata_int[7]),.T2I1(NET_44_CAND4_BLSBR_12_tpGCLKBUF),.T2I2(NET_45),.T2I3(m1_oper1_rdata_int[7]),.TB2S(GND),.C2Z(NET_474),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_L31_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m1_oper1_rdata_int[0]),.T3I1(m1_oper0_rdata_int[0]),.T3I2(NET_45),.T3I3(NET_44_CAND4_BLSBR_12_tpGCLKBUF),.C3Z(NET_116),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L32_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_43_CAND3_BLSBR_12_tpGCLKBUF),.B0I1(m1_oper0_rdata_int[18]),.B0I2(m1_coef_rdata_int[18]),.B0I3(NET_45),.T0I0(NET_44_CAND4_BLSBR_12_tpGCLKBUF),.T0I1(m1_oper0_rdata_int[6]),.T0I2(NET_45),.T0I3(m1_oper1_rdata_int[6]),.TB0S(GND),.B0Z(NET_364),.C0Z(NET_640),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_L32_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m1_coef_rdata_int[21]),.T1I1(m1_oper0_rdata_int[21]),.T1I2(NET_43_CAND3_BLSBR_12_tpGCLKBUF),.T1I3(NET_45),.C1Z(NET_419),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_L32_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_oper0_rdata_int[23]),.B2I1(NET_45),.B2I2(NET_43_CAND3_BLSBR_12_tpGCLKBUF),.B2I3(m1_coef_rdata_int[23]),.T2I0(m1_oper1_rdata_int[12]),.T2I1(NET_44_CAND4_BLSBR_12_tpGCLKBUF),.T2I2(m1_oper0_rdata_int[12]),.T2I3(NET_45),.TB2S(GND),.B2Z(NET_455),.C2Z(NET_228),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_L32_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m1_oper0_rdata_int[17]),.T3I1(m1_coef_rdata_int[17]),.T3I2(NET_43_CAND3_BLSBR_12_tpGCLKBUF),.T3I3(NET_45),.C3Z(NET_346),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M1_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.B0I1(NET_41),.B0I2(m0_coef_rdata_int[28]),.B0I3(m0_oper1_rdata_int[28]),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(m0_oper1_rdata_int[23]),.T0I1(m0_coef_rdata_int[23]),.T0I2(NET_41),.T0I3(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.TB0S(GND),.B0Z(NET_566),.C0Z(NET_457),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M1_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.T1I0(m0_coef_rdata_int[31]),.T1I1(m0_oper1_rdata_int[31]),.T1I2(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.T1I3(NET_41),.C1Z(NET_615),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_M1_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.T2I0(m0_oper1_rdata_int[26]),.T2I1(m0_coef_rdata_int[26]),.T2I2(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.T2I3(NET_41),.TB2S(GND),.C2Z(NET_531),.Q2Z(m0_coef_wdata_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_M1_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.T3I1(NET_41),.T3I2(m0_oper1_rdata_int[22]),.T3I3(m0_coef_rdata_int[22]),.C3Z(NET_439),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M3_0 (.tFragBitInfo(16'b0010101000000000),.bFragBitInfo(16'b0100110000000000),.B0I0(NET_41),.B0I1(NET_39),.B0I2(m0_coef_rdata_int[1]),.B0I3(NET_40),.T0I0(NET_658),.T0I1(NET_41),.T0I2(m0_coef_rdata_int[5]),.T0I3(NET_657),.TB0S(GND),.B0Z(NET_42),.C0Z(NET_659),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_M3_1 (.tFragBitInfo(16'b1010101011111111),.bFragBitInfo(16'b1111001110100011),.B1I0(lint_ADDR_int_13__CAND4_TLSTR_13_tpGCLKBUF),.B1I1(lint_ADDR_int[11]),.B1I2(apb_fsm[0]),.B1I3(lint_ADDR_int_14__CAND5_TLSTR_13_tpGCLKBUF),.T1I0(apb_fsm[0]),.T1I1(lint_ADDR_int_14__CAND5_TLSTR_13_tpGCLKBUF),.T1I2(lint_ADDR_int_13__CAND4_TLSTR_13_tpGCLKBUF),.T1I3(lint_ADDR_int[11]),.TB1S(m0_oper0_rdata_int[1]),.C1Z(NET_47),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_M3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_45),.B2I1(m1_oper0_rdata_int[5]),.B2I2(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.B2I3(m0_oper1_rdata_int[5]),.T2I0(NET_45),.T2I1(m1_oper0_rdata_int[5]),.T2I2(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.T2I3(m0_oper1_rdata_int[5]),.TB2S(NET_660),.C2Z(NET_658),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_M3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.B3I1(m1_oper0_rdata_int[1]),.B3I2(m0_oper1_rdata_int[1]),.B3I3(NET_45),.T3I0(m0_oper1_rdata_int[1]),.T3I1(NET_45),.T3I2(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.T3I3(m1_oper0_rdata_int[1]),.TB3S(NET_47),.C3Z(NET_40),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_M4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_oper0_rdata_int[11]),.B2I1(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.B2I2(NET_45),.B2I3(m0_oper1_rdata_int[11]),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.T2I0(m1_oper0_rdata_int[11]),.T2I1(NET_46_CAND1_TLSTR_13_tpGCLKBUF),.T2I2(NET_45),.T2I3(m0_oper1_rdata_int[11]),.TB2S(NET_206),.C2Z(NET_204),.Q2Z(m0_coef_wdata_dup_0[31]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_M4_3 (.tFragBitInfo(16'b0010000010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_204),.T3I1(m0_coef_rdata_int[11]),.T3I2(NET_203),.T3I3(NET_41),.C3Z(NET_205),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M5_0 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0111000000000000),.B0I0(m0_coef_rdata_int[3]),.B0I1(NET_41),.B0I2(NET_697),.B0I3(NET_696),.T0I0(apb_fsm[0]),.T0I1(GND),.T0I2(lint_ADDR_int_13__CAND4_TLSTR_13_tpGCLKBUF),.T0I3(lint_ADDR_int[12]),.TB0S(GND),.B0Z(NET_698),.C0Z(NET_41),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_M5_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[12]),.T1I1(NET_144),.T1I2(lint_ADDR_int_13__CAND4_TLSTR_13_tpGCLKBUF),.T1I3(NET_65),.C1Z(nx15998z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_M5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M5_3 (.tFragBitInfo(16'b0000100010001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_678),.T3I1(NET_677),.T3I2(m0_coef_rdata_int[4]),.T3I3(NET_41),.C3Z(NET_679),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M7_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B0I0(m0_m1_outsel_dup_0[4]),.B0I1(NET_62),.B0I2(tcdm_rdata_p0_int[4]),.B0I3(NET_63),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p0_int[8]),.T0I1(NET_62),.T0I2(m0_m1_control[8]),.T0I3(NET_63),.TB0S(GND),.B0Z(NET_682),.C0Z(NET_288),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[9]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_control[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_control[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M7_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[4]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_62),.T3I1(tcdm_rdata_p0_int[9]),.T3I2(m0_m1_control[9]),.T3I3(NET_63),.TB3S(GND),.C3Z(NET_167),.Q3Z(tcdm_result_p0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_outsel_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_63),.B2I1(tcdm_rdata_p0_int[10]),.B2I2(NET_62),.B2I3(m0_m1_control[10]),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.B2Z(NET_189),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_control[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M9_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B0I0(m0_coef_rdata_int[2]),.B0I1(NET_41),.B0I2(NET_43),.B0I3(m1_coef_rdata_int[2]),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(m1_coef_rdata_int[6]),.T0I1(NET_41),.T0I2(NET_43),.T0I3(m0_coef_rdata_int[6]),.TB0S(GND),.B0Z(NET_720),.C0Z(NET_639),.Q0Z(m0_m1_control[11]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M9_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_63),.T1I1(m0_m1_control[11]),.T1I2(NET_62),.T1I3(tcdm_rdata_p0_int[11]),.C1Z(NET_208),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_M9_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B2I0(m0_coef_rdata_int[7]),.B2I1(m1_coef_rdata_int[7]),.B2I2(NET_43),.B2I3(NET_41),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(m1_coef_rdata_int[0]),.T2I1(m0_coef_rdata_int[0]),.T2I2(NET_43),.T2I3(NET_41),.TB2S(GND),.B2Z(NET_473),.C2Z(NET_115),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_M9_3 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_15_CAND5_TLSBR_13_tpGCLKBUF),.T3I1(GND),.T3I2(GND),.T3I3(NET_8),.C3Z(NET_62),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B1I0(apb_fsm[0]),.B1I1(lint_ADDR_int[8]),.B1I2(lint_ADDR_int[2]),.B1I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[2]),.T1I1(lint_ADDR_int[11]),.T1I2(apb_fsm[0]),.T1I3(lint_ADDR_int[8]),.TB1S(lint_ADDR_int[7]),.C1Z(NET_89),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_M10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[10]),.Q3EN(tcdm_valid_p0_int_CAND1_TLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M11_0 (.tFragBitInfo(16'b1010000000000000),.bFragBitInfo(16'b0010000000000000),.B0I0(NET_615),.B0I1(m0_oper0_rdata_int[31]),.B0I2(NET_754),.B0I3(NET_614),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[11]),.Q0EN(tcdm_valid_p0_int_CAND1_TLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_615),.T0I1(m0_oper0_rdata_int[31]),.T0I2(NET_754),.T0I3(NET_614),.TB0S(NET_117),.C0Z(NET_606),.Q0Z(tcdm_result_p0[11]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M11_1 (.tFragBitInfo(16'b1000100000000000),.bFragBitInfo(16'b0100000000000000),.B1I0(m0_oper0_rdata_int[16]),.B1I1(NET_325),.B1I2(NET_324),.B1I3(NET_744),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[13]),.Q1EN(tcdm_valid_p0_int_CAND1_TLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_324),.T1I1(NET_744),.T1I2(m0_oper0_rdata_int[16]),.T1I3(NET_325),.TB1S(NET_117),.C1Z(NET_315),.Q1Z(tcdm_result_p0[13]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M11_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000010000),.B2I0(GND),.B2I1(lint_ADDR_int[13]),.B2I2(apb_fsm[0]),.B2I3(lint_ADDR_int[14]),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_10),.T2I1(GND),.T2I2(GND),.T2I3(NET_38),.TB2S(GND),.B2Z(NET_117),.C2Z(NET_63),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_M11_3 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_10),.T3I1(lint_ADDR_int[11]),.T3I2(GND),.T3I3(NET_38),.C3Z(NET_112),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M12_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_6),.T0I1(NET_36),.T0I2(m0_m0_control[20]),.T0I3(tcdm_rdata_p2_int[20]),.TB0S(GND),.C0Z(NET_403),.Q0Z(m0_m1_sat_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M12_1 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(NET_38),.T1I2(GND),.T1I3(NET_8),.C1Z(NET_36),.Q1Z(m0_m0_control[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_M12_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000100000000),.B2I0(lint_ADDR_int[3]),.B2I1(lint_ADDR_int[5]),.B2I2(lint_ADDR_int[6]),.B2I3(lint_ADDR_int[4]),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_401),.T2I1(NET_402),.T2I2(NET_400),.T2I3(NET_403),.TB2S(GND),.B2Z(NET_38),.C2Z(NET_388),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_M12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_mode_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M13_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(m0_m0_reset_dup_0),.B0I1(NET_6),.B0I2(tcdm_rdata_p2_int[31]),.B0I3(NET_36),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.T0I0(NET_617),.T0I1(NET_616),.T0I2(NET_619),.T0I3(NET_618),.TB0S(GND),.B0Z(NET_619),.C0Z(NET_604),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M13_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B1I0(NET_315),.B1I1(NET_312),.B1I2(NET_313),.B1I3(NET_314),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64_CAND2_TLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.T1I0(NET_313),.T1I1(NET_314),.T1I2(NET_315),.T1I3(NET_312),.TB1S(NET_316),.Q1Z(lint_RDATA_dup_0[16]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_M13_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_605),.B2I1(NET_603),.B2I2(NET_606),.B2I3(NET_604),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64_CAND2_TLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.T2I0(NET_605),.T2I1(NET_603),.T2I2(NET_606),.T2I3(NET_604),.TB2S(NET_607),.Q2Z(lint_RDATA_dup_0[31]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_M13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100010001000),.B0I0(NET_455),.B0I1(NET_456),.B0I2(NET_124_CAND4_TLSBR_13_tpGCLKBUF),.B0I3(tcdm_rdata_p0_int[23]),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_455),.T0I1(NET_456),.T0I2(NET_124_CAND4_TLSBR_13_tpGCLKBUF),.T0I3(tcdm_rdata_p0_int[23]),.TB0S(NET_457),.C0Z(NET_440),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_m0_tc_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M14_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000001000000),.B2I0(lint_ADDR_int[11]),.B2I1(NET_38),.B2I2(NET_8),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_rdata_int[23]),.T2I1(NET_117),.T2I2(NET_44),.T2I3(m0_oper0_rdata_int[23]),.TB2S(GND),.B2Z(NET_108),.C2Z(NET_456),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_M14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_reset_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000010100000),.B0I0(NET_438),.B0I1(NET_124_CAND4_TLSBR_13_tpGCLKBUF),.B0I2(NET_437),.B0I3(tcdm_rdata_p0_int[22]),.T0I0(NET_438),.T0I1(NET_124_CAND4_TLSBR_13_tpGCLKBUF),.T0I2(NET_437),.T0I3(tcdm_rdata_p0_int[22]),.TB0S(NET_439),.C0Z(NET_422),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_M15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000010100000),.B1I0(NET_365),.B1I1(NET_124_CAND4_TLSBR_13_tpGCLKBUF),.B1I2(NET_364),.B1I3(tcdm_rdata_p0_int[18]),.T1I0(NET_364),.T1I1(tcdm_rdata_p0_int[18]),.T1I2(NET_365),.T1I3(NET_124_CAND4_TLSBR_13_tpGCLKBUF),.TB1S(NET_366),.C1Z(NET_349),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_M15_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_oper1_rdata_int[22]),.B2I1(m0_oper0_rdata_int[22]),.B2I2(NET_44),.B2I3(NET_117),.T2I0(m0_oper0_rdata_int[28]),.T2I1(NET_44),.T2I2(m1_oper1_rdata_int[28]),.T2I3(NET_117),.TB2S(GND),.B2Z(NET_438),.C2Z(NET_565),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_M15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000010100000),.B3I0(NET_564),.B3I1(tcdm_rdata_p0_int[28]),.B3I2(NET_565),.B3I3(NET_124_CAND4_TLSBR_13_tpGCLKBUF),.T3I0(NET_565),.T3I1(NET_124_CAND4_TLSBR_13_tpGCLKBUF),.T3I2(NET_564),.T3I3(tcdm_rdata_p0_int[28]),.TB3S(NET_566),.C3Z(NET_549),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_M16_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_109),.B0I1(NET_108),.B0I2(tcdm_rdata_p2_int[0]),.B0I3(m0_m0_outsel_dup_0[0]),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p2_int[18]),.T0I1(m0_m1_sat_dup_0),.T0I2(NET_112),.T0I3(NET_109),.TB0S(GND),.B0Z(NET_106),.C0Z(NET_360),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M16_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[17]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p2_int[19]),.T1I1(m0_m1_control[19]),.T1I2(NET_112),.T1I3(NET_109),.TB1S(GND),.C1Z(NET_379),.Q1Z(tcdm_result_p2[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M16_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B2I0(tcdm_rdata_p2_int[12]),.B2I1(NET_108),.B2I2(m0_m0_mode_dup_0[0]),.B2I3(NET_109),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_109),.T2I1(m0_m1_clr_dup_0),.T2I2(NET_112),.T2I3(tcdm_rdata_p2_int[17]),.TB2S(GND),.B2Z(NET_223),.C2Z(NET_342),.Q2Z(m0_m1_control[19]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_M16_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p2_int[6]),.T3I1(NET_108),.T3I2(m0_m0_tc_dup_0),.T3I3(NET_109),.C3Z(NET_635),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M17_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[28]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_112),.T0I1(NET_109),.T0I2(tcdm_rdata_p2_int[28]),.T0I3(m0_m1_control[28]),.TB0S(GND),.C0Z(NET_560),.Q0Z(m0_m1_control[28]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_109),.B2I1(NET_108),.B2I2(m0_m0_outsel_dup_0[2]),.B2I3(tcdm_rdata_p2_int[2]),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[26]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B2Z(NET_716),.Q2Z(tcdm_result_p2[26]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B3I0(tcdm_result_p2[26]),.B3I1(NET_82),.B3I2(m0_m0_dataout_int[26]),.B3I3(NET_334),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx19726z1_CAND2_BLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_dataout_int[26]),.T3I1(NET_334),.T3I2(tcdm_result_p2[26]),.T3I3(NET_82),.TB3S(NET_518),.C3Z(NET_516),.Q3Z(m0_coef_wmode_dup_0[1]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M18_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_112),.B0I1(NET_109),.B0I2(m0_m1_control[23]),.B0I3(tcdm_rdata_p2_int[23]),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[23]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p2_int[24]),.T0I1(NET_112),.T0I2(m0_m1_control[24]),.T0I3(NET_109),.TB0S(GND),.B0Z(NET_451),.C0Z(NET_490),.Q0Z(tcdm_result_p2[23]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_control[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_82),.B2I1(tcdm_result_p2[28]),.B2I2(m0_m0_dataout_int[28]),.B2I3(NET_334),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[28]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_82),.T2I1(tcdm_result_p2[28]),.T2I2(m0_m0_dataout_int[28]),.T2I3(NET_334),.TB2S(NET_553),.C2Z(NET_551),.Q2Z(tcdm_result_p2[28]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_M18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B3I0(m0_m0_dataout_int[23]),.B3I1(NET_334),.B3I2(tcdm_result_p2[23]),.B3I3(NET_82),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p2[23]),.T3I1(NET_82),.T3I2(m0_m0_dataout_int[23]),.T3I3(NET_334),.TB3S(NET_444),.C3Z(NET_442),.Q3Z(m0_m1_control[23]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_65),.B0I1(NET_68),.B0I2(NET_66),.B0I3(lint_ADDR_int[3]),.T0I0(NET_65),.T0I1(NET_68),.T0I2(NET_66),.T0I3(lint_ADDR_int[3]),.TB0S(lint_ADDR_int[4]),.C0Z(nx28356z1),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_M19_1 (.tFragBitInfo(16'b1111101011111010),.bFragBitInfo(16'b1111100011111010),.B1I0(NET_726),.B1I1(NET_66),.B1I2(NET_622),.B1I3(NET_755),.T1I0(NET_622),.T1I1(NET_755),.T1I2(NET_726),.T1I3(NET_66),.TB1S(NET_620),.C1Z(nx49808z64),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_M19_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000010000),.B2I0(GND),.B2I1(GND),.B2I2(apb_fsm[1]),.B2I3(apb_fsm[0]),.T2I0(lint_ADDR_int[0]),.T2I1(lint_ADDR_int[1]),.T2I2(GND),.T2I3(lint_ADDR_int[9]),.TB2S(GND),.B2Z(NET_726),.C2Z(NET_71),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_M19_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_7),.T3I1(lint_ADDR_int[7]),.T3I2(lint_ADDR_int[2]),.T3I3(NET_19),.C3Z(NET_33),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M20_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0010001000000011),.B0I0(lint_ADDR_int[14]),.B0I1(GND),.B0I2(lint_ADDR_int[12]),.B0I3(lint_ADDR_int[13]),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_505),.T0I1(NET_502),.T0I2(NET_503),.T0I3(NET_504),.TB0S(GND),.B0Z(NET_621),.C0Z(NET_499),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_537),.B2I1(NET_539),.B2I2(NET_538),.B2I3(NET_540),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B2Z(NET_534),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M20_3 (.tFragBitInfo(16'b1000100000000000),.bFragBitInfo(16'b1100000001000000),.B3I0(NET_621),.B3I1(apb_fsm[1]),.B3I2(apb_fsm[0]),.B3I3(NET_171),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(apb_fsm[0]),.T3I1(NET_171),.T3I2(NET_621),.T3I3(apb_fsm[1]),.TB3S(NET_141),.C3Z(NET_622),.Q3Z(m1_m1_mode_dup_0[0]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_611),.B0I1(NET_610),.B0I2(NET_609),.B0I3(NET_608),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B0Z(NET_605),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M21_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_590),.T1I1(NET_591),.T1I2(NET_593),.T1I3(NET_592),.TB1S(GND),.C1Z(NET_587),.Q1Z(m1_m1_tc_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_sat_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M22_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.B0I0(NET_17_CAND3_BLSTR_13_tpGCLKBUF),.B0I1(NET_28_CAND4_BLSTR_13_tpGCLKBUF),.B0I2(m1_m1_control[20]),.B0I3(m1_ram_control[20]),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_17_CAND3_BLSTR_13_tpGCLKBUF),.T0I1(NET_28_CAND4_BLSTR_13_tpGCLKBUF),.T0I2(m1_m1_control[20]),.T0I3(m1_ram_control[20]),.TB0S(NET_396),.C0Z(NET_394),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_control[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx19726z1_CAND2_BLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_rmode_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M22_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[20]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_394),.T3I1(NET_393),.T3I2(NET_395),.T3I3(NET_392),.TB3S(GND),.C3Z(NET_389),.Q3Z(m1_ram_control[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_control[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M25_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_control[27]),.T3I1(NET_33),.T3I2(m1_m1_dataout_int[27]),.T3I3(NET_32_CAND5_BLSBR_13_tpGCLKBUF),.C3Z(NET_538),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M26_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(m1_m1_dataout_int[20]),.T0I1(NET_32_CAND5_BLSBR_13_tpGCLKBUF),.T0I2(m1_m0_control[20]),.T0I3(NET_33),.TB0S(GND),.C0Z(NET_393),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_control[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M27_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(m1_m1_dataout_int[25]),.T0I1(NET_32_CAND5_BLSBR_13_tpGCLKBUF),.T0I2(m1_m0_control[25]),.T0I3(NET_33),.TB0S(GND),.C0Z(NET_503),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_control[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M28_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_65),.T1I1(GND),.T1I2(NET_171),.T1I3(lint_ADDR_int[13]),.TB1S(GND),.C1Z(nx33579z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_M28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M29_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_dataout_int[30]),.T1I1(NET_33),.T1I2(m1_m0_control[30]),.T1I3(NET_32_CAND5_BLSBR_13_tpGCLKBUF),.TB1S(GND),.C1Z(NET_591),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_M29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_control[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M29_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_32_CAND5_BLSBR_13_tpGCLKBUF),.T3I1(NET_33),.T3I2(m1_m0_control[10]),.T3I3(m1_m1_dataout_int[10]),.TB3S(GND),.C3Z(NET_182),.Q3Z(m1_m0_control[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_32_CAND5_BLSBR_13_tpGCLKBUF),.B0I1(NET_33),.B0I2(m1_m0_reset_dup_0),.B0I3(m1_m1_dataout_int[31]),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B0Z(NET_609),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M30_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_dataout_int[13]),.T1I1(NET_32_CAND5_BLSBR_13_tpGCLKBUF),.T1I2(m1_m0_mode_dup_0[1]),.T1I3(NET_33),.TB1S(GND),.C1Z(NET_241),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_M30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_reset_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(m1_m0_mode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.B0I1(m1_coef_rdata_int[13]),.B0I2(NET_44_CAND4_BLSBR_13_tpGCLKBUF),.B0I3(m1_oper1_rdata_int[13]),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B0Z(NET_243),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M31_1 (.tFragBitInfo(16'b1010101011111111),.bFragBitInfo(16'b1111001110100011),.B1I0(lint_ADDR_int[12]),.B1I1(lint_ADDR_int[11]),.B1I2(apb_fsm[0]),.B1I3(lint_ADDR_int[13]),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(apb_fsm[0]),.T1I1(lint_ADDR_int[13]),.T1I2(lint_ADDR_int[12]),.T1I3(lint_ADDR_int[11]),.TB1S(m1_oper0_rdata_int[27]),.C1Z(NET_749),.Q1Z(m1_coef_wdata_dup_0[31]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M31_2 (.tFragBitInfo(16'b1010101011111111),.bFragBitInfo(16'b1010100011111101),.B2I0(apb_fsm[0]),.B2I1(lint_ADDR_int[13]),.B2I2(lint_ADDR_int[12]),.B2I3(lint_ADDR_int[11]),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(apb_fsm[0]),.T2I1(lint_ADDR_int[13]),.T2I2(lint_ADDR_int[12]),.T2I3(lint_ADDR_int[11]),.TB2S(m1_oper0_rdata_int[25]),.C2Z(NET_747),.Q2Z(m1_coef_wdata_dup_0[13]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_M31_3 (.tFragBitInfo(16'b0010001010101010),.bFragBitInfo(16'b0001000001010000),.B3I0(m1_oper1_rdata_int[31]),.B3I1(m1_coef_rdata_int[31]),.B3I2(NET_753),.B3I3(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_753),.T3I1(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.T3I2(m1_oper1_rdata_int[31]),.T3I3(m1_coef_rdata_int[31]),.TB3S(NET_44_CAND4_BLSBR_13_tpGCLKBUF),.C3Z(NET_754),.Q3Z(m1_coef_wdata_dup_0[30]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(m1_oper1_rdata_int[9]),.B0I1(m1_coef_rdata_int[9]),.B0I2(NET_44_CAND4_BLSBR_13_tpGCLKBUF),.B0I3(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B0Z(NET_162),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M32_1 (.tFragBitInfo(16'b0111000001110000),.bFragBitInfo(16'b0000001000100010),.B1I0(NET_743),.B1I1(m1_oper1_rdata_int[16]),.B1I2(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.B1I3(m1_coef_rdata_int[16]),.CD1S(VCC),.Q1DI(lint_WDATA_int[26]),.Q1EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.T1I1(m1_coef_rdata_int[16]),.T1I2(NET_743),.T1I3(m1_oper1_rdata_int[16]),.TB1S(NET_44_CAND4_BLSBR_13_tpGCLKBUF),.C1Z(NET_744),.Q1Z(m1_coef_wdata_dup_0[26]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M32_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_oper0_rdata_int[19]),.B2I1(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.B2I2(NET_45),.B2I3(m1_coef_rdata_int[19]),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_rdata_int[8]),.T2I1(m1_coef_rdata_int[8]),.T2I2(NET_44_CAND4_BLSBR_13_tpGCLKBUF),.T2I3(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.TB2S(GND),.B2Z(NET_383),.C2Z(NET_283),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_M32_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(m1_coef_rdata_int[22]),.T3I1(NET_43_CAND3_BLSBR_13_tpGCLKBUF),.T3I2(m1_oper0_rdata_int[22]),.T3I3(NET_45),.TB3S(GND),.C3Z(NET_437),.Q3Z(m1_coef_wdata_dup_0[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_N1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[12]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N1_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(m0_oper1_rdata_int[17]),.T1I1(NET_41),.T1I2(m0_coef_rdata_int[17]),.T1I3(NET_46_CAND1_TLSTR_14_tpGCLKBUF),.TB1S(GND),.C1Z(NET_348),.Q1Z(m0_coef_wdata_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N1_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.T2I0(m0_coef_rdata_int[27]),.T2I1(NET_41),.T2I2(NET_46_CAND1_TLSTR_14_tpGCLKBUF),.T2I3(m0_oper1_rdata_int[27]),.TB2S(GND),.C2Z(NET_544),.Q2Z(m0_coef_wdata_dup_0[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[27]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[23]),.Q1EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[23]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[21]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000000000000),.B0I0(lint_ADDR_int_14__CAND5_TLSTR_14_tpGCLKBUF),.B0I1(lint_WEN_int),.B0I2(lint_ADDR_int_13__CAND4_TLSTR_14_tpGCLKBUF),.B0I3(lint_ADDR_int[12]),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.B0Z(NET_311),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N5_1 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int_14__CAND5_TLSTR_14_tpGCLKBUF),.T1I1(lint_WEN_int),.T1I2(lint_ADDR_int_13__CAND4_TLSTR_14_tpGCLKBUF),.T1I3(lint_ADDR_int[12]),.TB1S(GND),.C1Z(NET_151),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_N5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_outsel_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_tc_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_csel_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N8_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p0_int[15]),.T1I1(m0_m1_csel_dup_0),.T1I2(NET_63),.T1I3(NET_62),.TB1S(GND),.C1Z(NET_307),.Q1Z(m0_m1_mode_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[14]),.Q0EN(tcdm_valid_p0_int_CAND1_TLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[15]),.Q1EN(tcdm_valid_p0_int_CAND1_TLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N10_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[13]),.T2I1(lint_ADDR_int[14]),.T2I2(apb_fsm[0]),.T2I3(GND),.TB2S(GND),.C2Z(NET_43),.Q2Z(m0_m0_outsel_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N11_0 (.tFragBitInfo(16'b1000100000000000),.bFragBitInfo(16'b0000100000000000),.B0I0(NET_398),.B0I1(NET_399),.B0I2(m0_oper0_rdata_int[20]),.B0I3(NET_746),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_398),.T0I1(NET_399),.T0I2(m0_oper0_rdata_int[20]),.T0I3(NET_746),.TB0S(NET_117),.C0Z(NET_390),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N11_1 (.tFragBitInfo(16'b1000000010000000),.bFragBitInfo(16'b0010000000000000),.B1I0(NET_597),.B1I1(m0_oper0_rdata_int[30]),.B1I2(NET_596),.B1I3(NET_752),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_596),.T1I1(NET_752),.T1I2(NET_597),.T1I3(m0_oper0_rdata_int[30]),.TB1S(NET_117),.C1Z(NET_588),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_N11_2 (.tFragBitInfo(16'b1100000000000000),.bFragBitInfo(16'b0100000000000000),.B2I0(m0_oper0_rdata_int[25]),.B2I1(NET_748),.B2I2(NET_508),.B2I3(NET_509),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(m0_oper0_rdata_int[25]),.T2I1(NET_748),.T2I2(NET_508),.T2I3(NET_509),.TB2S(NET_117),.C2Z(NET_500),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_N11_3 (.tFragBitInfo(16'b1010000000000000),.bFragBitInfo(16'b0000000010000000),.B3I0(NET_543),.B3I1(NET_544),.B3I2(NET_750),.B3I3(m0_oper0_rdata_int[27]),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(NET_750),.T3I1(m0_oper0_rdata_int[27]),.T3I2(NET_543),.T3I3(NET_544),.TB3S(NET_117),.C3Z(NET_535),.Q3Z(m0_m0_control[25]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_N12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_510),.B0I1(NET_511),.B0I2(NET_513),.B0I3(NET_512),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.B0Z(NET_498),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N12_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B1I0(NET_387),.B1I1(NET_388),.B1I2(NET_389),.B1I3(NET_390),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64_CAND2_TLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.T1I0(NET_389),.T1I1(NET_390),.T1I2(NET_387),.T1I3(NET_388),.TB1S(NET_391),.Q1Z(lint_RDATA_dup_0[20]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_N12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_36),.B2I1(m0_m0_control[25]),.B2I2(NET_6),.B2I3(tcdm_rdata_p2_int[25]),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.B2Z(NET_513),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N12_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_499),.B3I1(NET_497),.B3I2(NET_500),.B3I3(NET_498),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z64_CAND2_TLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.T3I0(NET_500),.T3I1(NET_498),.T3I2(NET_499),.T3I3(NET_497),.TB3S(NET_501),.Q3Z(lint_RDATA_dup_0[25]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_N13_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.T0I0(NET_601),.T0I1(NET_599),.T0I2(NET_600),.T0I3(NET_598),.TB0S(GND),.C0Z(NET_586),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N13_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B1I0(NET_588),.B1I1(NET_586),.B1I2(NET_585),.B1I3(NET_587),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z64_CAND2_TLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.T1I0(NET_585),.T1I1(NET_587),.T1I2(NET_588),.T1I3(NET_586),.TB1S(NET_589),.Q1Z(lint_RDATA_dup_0[30]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_N13_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_535),.B2I1(NET_534),.B2I2(NET_533),.B2I3(NET_532),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z64_CAND2_TLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.T2I0(NET_535),.T2I1(NET_534),.T2I2(NET_533),.T2I3(NET_532),.TB2S(NET_536),.Q2Z(lint_RDATA_dup_0[27]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_N13_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.T3I0(NET_548),.T3I1(NET_545),.T3I2(NET_547),.T3I3(NET_546),.TB3S(GND),.C3Z(NET_533),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_N14_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p2_int[30]),.T0I1(NET_6),.T0I2(NET_36),.T0I3(m0_m0_control[30]),.TB0S(GND),.C0Z(NET_601),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0111000000000000),.B1I0(tcdm_rdata_p0_int[24]),.B1I1(NET_124_CAND4_TLSBR_14_tpGCLKBUF),.B1I2(NET_495),.B1I3(NET_494),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_495),.T1I1(NET_494),.T1I2(tcdm_rdata_p0_int[24]),.T1I3(NET_124_CAND4_TLSBR_14_tpGCLKBUF),.TB1S(NET_496),.C1Z(NET_479),.Q1Z(m0_m0_control[30]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N14_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B2I0(m0_oper0_rdata_int[24]),.B2I1(m1_oper1_rdata_int[24]),.B2I2(NET_117),.B2I3(NET_44),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(m0_m0_control[27]),.T2I1(NET_6),.T2I2(tcdm_rdata_p2_int[27]),.T2I3(NET_36),.TB2S(GND),.B2Z(NET_495),.C2Z(NET_548),.Q2Z(m0_m0_control[27]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_N14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N15_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B0I0(m1_oper1_rdata_int[19]),.B0I1(NET_44),.B0I2(m0_oper0_rdata_int[19]),.B0I3(NET_117),.T0I0(m1_oper1_rdata_int[18]),.T0I1(NET_44),.T0I2(m0_oper0_rdata_int[18]),.T0I3(NET_117),.TB0S(GND),.B0Z(NET_384),.C0Z(NET_365),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_N15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0111000000000000),.B1I0(NET_124_CAND4_TLSBR_14_tpGCLKBUF),.B1I1(tcdm_rdata_p0_int[17]),.B1I2(NET_347),.B1I3(NET_346),.T1I0(NET_347),.T1I1(NET_346),.T1I2(NET_124_CAND4_TLSBR_14_tpGCLKBUF),.T1I3(tcdm_rdata_p0_int[17]),.TB1S(NET_348),.C1Z(NET_330),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_N15_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000100000000000),.B2I0(tcdm_rdata_p1_int[25]),.B2I1(NET_15_CAND5_TLSBR_14_tpGCLKBUF),.B2I2(GND),.B2I3(NET_10),.T2I0(m0_oper0_rdata_int[17]),.T2I1(NET_44),.T2I2(NET_117),.T2I3(m1_oper1_rdata_int[17]),.TB2S(GND),.B2Z(NET_506),.C2Z(NET_347),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_N15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010101000000000),.B3I0(NET_383),.B3I1(tcdm_rdata_p0_int[19]),.B3I2(NET_124_CAND4_TLSBR_14_tpGCLKBUF),.B3I3(NET_384),.T3I0(NET_124_CAND4_TLSBR_14_tpGCLKBUF),.T3I1(NET_384),.T3I2(NET_383),.T3I3(tcdm_rdata_p0_int[19]),.TB3S(NET_385),.C3Z(NET_368),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_N16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_96),.B0I1(tcdm_result_p3[17]),.B0I2(NET_99),.B0I3(fpgaio_out_dup_0[49]),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_96),.T0I1(tcdm_result_p3[17]),.T0I2(NET_99),.T0I3(fpgaio_out_dup_0[49]),.TB0S(NET_339),.C0Z(NET_336),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B1I0(NET_99),.B1I1(fpgaio_out_dup_0[50]),.B1I2(NET_96),.B1I3(tcdm_result_p3[18]),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[18]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_96),.T1I1(tcdm_result_p3[18]),.T1I2(NET_99),.T1I3(fpgaio_out_dup_0[50]),.TB1S(NET_357),.C1Z(NET_354),.Q1Z(tcdm_result_p2[18]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000010000000000),.B2I0(GND),.B2I1(NET_125),.B2I2(GND),.B2I3(NET_8),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.B2Z(NET_124),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_outsel_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001000000000000),.B0I0(GND),.B0I1(GND),.B0I2(NET_8),.B0I3(NET_110),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B0Z(NET_109),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N17_1 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[6]),.T1I1(NET_146),.T1I2(NET_135),.T1I3(lint_ADDR_int[5]),.TB1S(GND),.C1Z(nx19726z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_N17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_96),.B2I1(fpgaio_out_dup_0[61]),.B2I2(tcdm_result_p3[29]),.B2I3(NET_99),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_96),.T2I1(fpgaio_out_dup_0[61]),.T2I2(tcdm_result_p3[29]),.T2I3(NET_99),.TB2S(NET_575),.C2Z(NET_572),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_N17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B3I0(lint_ADDR_int[4]),.B3I1(lint_ADDR_int[5]),.B3I2(lint_ADDR_int[6]),.B3I3(lint_ADDR_int[11]),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx19726z1_CAND2_BLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[6]),.T3I1(lint_ADDR_int[11]),.T3I2(lint_ADDR_int[4]),.T3I3(lint_ADDR_int[5]),.TB3S(lint_ADDR_int[3]),.C3Z(NET_110),.Q3Z(m0_oper1_wmode_dup_0[1]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_N18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(tcdm_result_p3[23]),.B0I1(fpgaio_out_dup_0[55]),.B0I2(NET_96),.B0I3(NET_99),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p3[23]),.T0I1(fpgaio_out_dup_0[55]),.T0I2(NET_96),.T0I3(NET_99),.TB0S(NET_448),.C0Z(NET_445),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B1I0(NET_96),.B1I1(NET_99),.B1I2(tcdm_result_p3[24]),.B1I3(fpgaio_out_dup_0[56]),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx19726z1_CAND2_BLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p3[24]),.T1I1(fpgaio_out_dup_0[56]),.T1I2(NET_96),.T1I3(NET_99),.TB1S(NET_487),.C1Z(NET_484),.Q1Z(m0_coef_wmode_dup_0[0]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N18_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_67),.B2I1(NET_66),.B2I2(GND),.B2I3(NET_145),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_67),.T2I1(NET_66),.T2I2(NET_68),.T2I3(NET_65),.TB2S(GND),.B2Z(nx40728z1),.C2Z(nx10775z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_N18_3 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_8),.T3I2(NET_7),.T3I3(GND),.TB3S(GND),.C3Z(NET_6),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_N19_0 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000000000010000),.B0I0(GND),.B0I1(lint_ADDR_int[3]),.B0I2(NET_75),.B0I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_133),.T0I1(NET_623),.T0I2(GND),.T0I3(NET_69),.TB0S(GND),.B0Z(NET_70),.C0Z(nx60509z1),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N19_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[4]),.T1I1(NET_134),.T1I2(NET_65),.T1I3(NET_66),.TB1S(GND),.C1Z(nx23147z1),.Q1Z(m1_m1_clr_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N19_2 (.tFragBitInfo(16'b0000000100001111),.bFragBitInfo(16'b0000000000001111),.B2I0(NET_62),.B2I1(NET_70),.B2I2(NET_147),.B2I3(NET_69),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx19726z1_CAND2_BLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_62),.T2I1(NET_70),.T2I2(NET_147),.T2I3(NET_69),.TB2S(NET_623),.C2Z(NET_755),.Q2Z(m0_coef_wdsel_dup_0),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N20_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.B0I0(NET_17_CAND3_BLSTR_14_tpGCLKBUF),.B0I1(m1_ram_control[27]),.B0I2(NET_28_CAND4_BLSTR_14_tpGCLKBUF),.B0I3(m1_m1_control[27]),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_17_CAND3_BLSTR_14_tpGCLKBUF),.T0I1(m1_ram_control[27]),.T0I2(NET_28_CAND4_BLSTR_14_tpGCLKBUF),.T0I3(m1_m1_control[27]),.TB0S(NET_541),.C0Z(NET_539),.Q0Z(m1_ram_control[27]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000010000),.B1I0(lint_ADDR_int[4]),.B1I1(lint_ADDR_int[7]),.B1I2(lint_ADDR_int[6]),.B1I3(lint_ADDR_int[11]),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[6]),.T1I1(lint_ADDR_int[11]),.T1I2(lint_ADDR_int[4]),.T1I3(lint_ADDR_int[7]),.TB1S(lint_ADDR_int[5]),.C1Z(NET_623),.Q1Z(m1_m1_control[25]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N20_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.B2I0(NET_17_CAND3_BLSTR_14_tpGCLKBUF),.B2I1(m1_ram_control[25]),.B2I2(NET_28_CAND4_BLSTR_14_tpGCLKBUF),.B2I3(m1_m1_control[25]),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_17_CAND3_BLSTR_14_tpGCLKBUF),.T2I1(m1_ram_control[25]),.T2I2(NET_28_CAND4_BLSTR_14_tpGCLKBUF),.T2I3(m1_m1_control[25]),.TB2S(NET_506),.C2Z(NET_504),.Q2Z(m1_ram_control[25]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_control[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N21_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.B0I0(NET_17_CAND3_BLSTR_14_tpGCLKBUF),.B0I1(NET_28_CAND4_BLSTR_14_tpGCLKBUF),.B0I2(m1_ram_control[31]),.B0I3(m1_m1_reset_dup_0),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_17_CAND3_BLSTR_14_tpGCLKBUF),.T0I1(NET_28_CAND4_BLSTR_14_tpGCLKBUF),.T0I2(m1_ram_control[31]),.T0I3(m1_m1_reset_dup_0),.TB0S(NET_612),.C0Z(NET_610),.Q0Z(m1_m1_control[30]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N21_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(apb_fsm[0]),.T1I1(lint_ADDR_int[12]),.T1I2(GND),.T1I3(lint_ADDR_int[14]),.C1Z(NET_44),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_N21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m1_ram_control[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N21_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.B3I0(m1_ram_control[30]),.B3I1(m1_m1_control[30]),.B3I2(NET_17_CAND3_BLSTR_14_tpGCLKBUF),.B3I3(NET_28_CAND4_BLSTR_14_tpGCLKBUF),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T3I0(NET_17_CAND3_BLSTR_14_tpGCLKBUF),.T3I1(NET_28_CAND4_BLSTR_14_tpGCLKBUF),.T3I2(m1_ram_control[30]),.T3I3(m1_m1_control[30]),.TB3S(NET_594),.C3Z(NET_592),.Q3Z(m1_ram_control[30]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_N22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m1_ram_control[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N22_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.B1I0(m1_m1_rnd_dup_0),.B1I1(NET_28_CAND4_BLSTR_14_tpGCLKBUF),.B1I2(m1_ram_control[16]),.B1I3(NET_17_CAND3_BLSTR_14_tpGCLKBUF),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(m1_ram_control[16]),.T1I1(NET_17_CAND3_BLSTR_14_tpGCLKBUF),.T1I2(m1_m1_rnd_dup_0),.T1I3(NET_28_CAND4_BLSTR_14_tpGCLKBUF),.TB1S(NET_321),.C1Z(NET_319),.Q1Z(m1_m1_reset_dup_0),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m1_m1_mode_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_rnd_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N23_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[12]),.T1I1(lint_ADDR_int[14]),.T1I2(lint_WEN_int),.T1I3(lint_ADDR_int[13]),.TB1S(GND),.C1Z(NET_646),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_N23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000000000000),.B2I0(lint_ADDR_int[12]),.B2I1(lint_ADDR_int[14]),.B2I2(lint_WEN_int),.B2I3(lint_ADDR_int[13]),.B2Z(NET_140),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N31_0 (.tFragBitInfo(16'b0111000001110000),.bFragBitInfo(16'b0000000001110000),.B0I0(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.B0I1(m1_coef_rdata_int[27]),.B0I2(NET_749),.B0I3(m1_oper1_rdata_int[27]),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.T0I1(m1_coef_rdata_int[27]),.T0I2(NET_749),.T0I3(m1_oper1_rdata_int[27]),.TB0S(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.C0Z(NET_750),.Q0Z(m1_coef_wdata_dup_0[29]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N31_1 (.tFragBitInfo(16'b0011111100000000),.bFragBitInfo(16'b0000010000001100),.B1I0(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.B1I1(NET_751),.B1I2(m1_oper1_rdata_int[30]),.B1I3(m1_coef_rdata_int[30]),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(m1_oper1_rdata_int[30]),.T1I1(m1_coef_rdata_int[30]),.T1I2(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.T1I3(NET_751),.TB1S(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.C1Z(NET_752),.Q1Z(m1_coef_wdata_dup_0[20]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N31_2 (.tFragBitInfo(16'b0000101010101010),.bFragBitInfo(16'b0000001000100010),.B2I0(NET_745),.B2I1(m1_oper1_rdata_int[20]),.B2I2(m1_coef_rdata_int[20]),.B2I3(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_745),.T2I1(m1_oper1_rdata_int[20]),.T2I2(m1_coef_rdata_int[20]),.T2I3(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.TB2S(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.C2Z(NET_746),.Q2Z(m1_coef_wdata_dup_0[21]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N32_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[28]),.Q0EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.T0I1(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.T0I2(m1_oper1_rdata_int[4]),.T0I3(m1_coef_rdata_int[4]),.TB0S(GND),.C0Z(NET_677),.Q0Z(m1_coef_wdata_dup_0[28]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N32_1 (.tFragBitInfo(16'b0101000011110000),.bFragBitInfo(16'b0000000000101010),.B1I0(NET_747),.B1I1(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.B1I2(m1_coef_rdata_int[25]),.B1I3(m1_oper1_rdata_int[25]),.CD1S(VCC),.Q1DI(lint_WDATA_int[23]),.Q1EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(m1_coef_rdata_int[25]),.T1I1(m1_oper1_rdata_int[25]),.T1I2(NET_747),.T1I3(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.TB1S(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.C1Z(NET_748),.Q1Z(m1_coef_wdata_dup_0[23]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_N32_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(m1_coef_rdata_int[1]),.T2I1(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.T2I2(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.T2I3(m1_oper1_rdata_int[1]),.TB2S(GND),.C2Z(NET_39),.Q2Z(m1_coef_wdata_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N32_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(m1_coef_rdata_int[3]),.T3I1(m1_oper1_rdata_int[3]),.T3I2(NET_43_CAND3_BLSBR_14_tpGCLKBUF),.T3I3(NET_44_CAND4_BLSBR_14_tpGCLKBUF),.TB3S(GND),.C3Z(NET_696),.Q3Z(m1_coef_wdata_dup_0[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_O1_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[0]),.Q0EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.T0I0(m0_oper1_rdata_int[30]),.T0I1(m0_coef_rdata_int[30]),.T0I2(NET_46_CAND1_TLSTR_15_tpGCLKBUF),.T0I3(NET_41),.TB0S(GND),.C0Z(NET_597),.Q0Z(m0_coef_waddr_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O1_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.T1I0(m0_oper1_rdata_int[21]),.T1I1(NET_41),.T1I2(m0_coef_rdata_int[21]),.T1I3(NET_46_CAND1_TLSTR_15_tpGCLKBUF),.TB1S(GND),.C1Z(NET_421),.Q1Z(m0_coef_wdata_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_O1_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_41),.T2I1(m0_coef_rdata_int[24]),.T2I2(NET_46_CAND1_TLSTR_15_tpGCLKBUF),.T2I3(m0_oper1_rdata_int[24]),.TB2S(GND),.C2Z(NET_496),.Q2Z(m0_coef_wdata_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[6]),.Q3EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_waddr_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000000000000),.B0I0(GND),.B0I1(NET_149),.B0I2(NET_65),.B0I3(lint_ADDR_int_13__CAND4_TLSTR_15_tpGCLKBUF),.B0Z(nx25587z1),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O5_2 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_311),.T2I1(GND),.T2I2(NET_142),.T2I3(NET_141),.TB2S(GND),.C2Z(nx32231z1),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_O5_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_151),.T3I1(GND),.T3I2(NET_142),.T3I3(NET_141),.C3Z(nx18281z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q0Z(m0_m1_osel_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_mode_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_63),.B0I1(NET_62),.B0I2(tcdm_rdata_p0_int[13]),.B0I3(m0_m1_mode_dup_0[1]),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.B0Z(NET_248),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O7_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.T1I0(NET_63),.T1I1(NET_62),.T1I2(tcdm_rdata_p0_int[5]),.T1I3(m0_m1_outsel_dup_0[5]),.TB1S(GND),.C1Z(NET_662),.Q1Z(m0_m1_outsel_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_O7_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_63),.B2I1(NET_62),.B2I2(tcdm_rdata_p0_int[3]),.B2I3(m0_m1_outsel_dup_0[3]),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_63),.T2I1(NET_62),.T2I2(m0_m1_outsel_dup_0[1]),.T2I3(tcdm_rdata_p0_int[1]),.TB2S(GND),.B2Z(NET_701),.C2Z(NET_54),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_O7_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_63),.T3I1(tcdm_rdata_p0_int[14]),.T3I2(m0_m1_osel_dup_0),.T3I3(NET_62),.C3Z(NET_268),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[5]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[1]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_63),.B0I1(NET_51),.B0I2(m0_m1_control[30]),.B0I3(tcdm_result_p3[30]),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.B0Z(NET_596),.Q0Z(m0_m1_control[27]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_control[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O11_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_63),.T2I1(NET_51),.T2I2(m0_m1_control[25]),.T2I3(tcdm_result_p3[25]),.TB2S(GND),.C2Z(NET_508),.Q2Z(m0_m1_control[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O11_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_63),.T3I1(NET_51),.T3I2(tcdm_result_p3[27]),.T3I3(m0_m1_control[27]),.C3Z(NET_543),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000000000000),.B0I0(NET_10),.B0I1(GND),.B0I2(tcdm_rdata_p1_int[20]),.B0I3(NET_15_CAND5_TLSBR_15_tpGCLKBUF),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[25]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.B0Z(NET_396),.Q0Z(tcdm_result_p1[25]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[30]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p3[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O12_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[25]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p0_int[20]),.T2I1(NET_50),.T2I2(NET_62),.T2I3(tcdm_result_p1[20]),.TB2S(GND),.C2Z(NET_391),.Q2Z(tcdm_result_p3[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O12_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[20]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p1[25]),.T3I1(NET_50),.T3I2(NET_62),.T3I3(tcdm_rdata_p0_int[25]),.C3Z(NET_501),.Q3Z(tcdm_result_p1[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O13_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[31]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(NET_62),.T0I1(tcdm_rdata_p0_int[31]),.T0I2(NET_50),.T0I3(tcdm_result_p1[31]),.TB0S(GND),.C0Z(NET_607),.Q0Z(tcdm_result_p1[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O13_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[30]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(NET_62),.T1I1(tcdm_result_p1[27]),.T1I2(tcdm_rdata_p0_int[27]),.T1I3(NET_50),.C1Z(NET_536),.Q1Z(tcdm_result_p1[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_62),.B2I1(tcdm_rdata_p0_int[30]),.B2I2(tcdm_result_p1[30]),.B2I3(NET_50),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[27]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.B2Z(NET_589),.Q2Z(tcdm_result_p1[27]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O13_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[16]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_62),.T3I1(tcdm_rdata_p0_int[16]),.T3I2(tcdm_result_p1[16]),.T3I3(NET_50),.TB3S(GND),.C3Z(NET_316),.Q3Z(tcdm_result_p1[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_O14_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(tcdm_result_p0[21]),.B0I1(NET_101),.B0I2(NET_89),.B0I3(tcdm_result_p1[21]),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[21]),.Q0EN(tcdm_valid_p0_int_CAND1_TLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p0[21]),.T0I1(NET_101),.T0I2(NET_89),.T0I3(tcdm_result_p1[21]),.TB0S(NET_15_CAND5_TLSBR_15_tpGCLKBUF),.C0Z(NET_412),.Q0Z(tcdm_result_p0[21]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O14_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B1I0(tcdm_result_p1[17]),.B1I1(tcdm_result_p0[17]),.B1I2(NET_89),.B1I3(NET_101),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[21]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(NET_89),.T1I1(NET_101),.T1I2(tcdm_result_p1[17]),.T1I3(tcdm_result_p0[17]),.TB1S(NET_15_CAND5_TLSBR_15_tpGCLKBUF),.C1Z(NET_339),.Q1Z(tcdm_result_p1[21]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_O14_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0100000000000000),.B2I0(GND),.B2I1(NET_15_CAND5_TLSBR_15_tpGCLKBUF),.B2I2(NET_10),.B2I3(tcdm_rdata_p1_int[16]),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[17]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p1_int[27]),.T2I1(NET_15_CAND5_TLSBR_15_tpGCLKBUF),.T2I2(GND),.T2I3(NET_10),.TB2S(GND),.B2Z(NET_321),.C2Z(NET_541),.Q2Z(tcdm_result_p1[17]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_O14_3 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[17]),.Q3EN(tcdm_valid_p0_int_CAND1_TLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p1_int[31]),.T3I1(NET_15_CAND5_TLSBR_15_tpGCLKBUF),.T3I2(GND),.T3I3(NET_10),.TB3S(GND),.C3Z(NET_612),.Q3Z(tcdm_result_p0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_O15_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_89),.B0I1(NET_101),.B0I2(tcdm_result_p1[29]),.B0I3(tcdm_result_p0[29]),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[29]),.Q0EN(tcdm_valid_p0_int_CAND1_TLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(NET_89),.T0I1(NET_101),.T0I2(tcdm_result_p1[29]),.T0I3(tcdm_result_p0[29]),.TB0S(NET_15_CAND5_TLSBR_15_tpGCLKBUF),.C0Z(NET_575),.Q0Z(tcdm_result_p0[29]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[29]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p1[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O15_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_101),.B2I1(NET_89),.B2I2(tcdm_result_p1[19]),.B2I3(tcdm_result_p0[19]),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[19]),.Q2EN(tcdm_valid_p0_int_CAND1_TLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_101),.T2I1(NET_89),.T2I2(tcdm_result_p1[19]),.T2I3(tcdm_result_p0[19]),.TB2S(NET_15_CAND5_TLSBR_15_tpGCLKBUF),.C2Z(NET_376),.Q2Z(tcdm_result_p0[19]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O15_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[19]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p1_int[30]),.T3I1(GND),.T3I2(NET_15_CAND5_TLSBR_15_tpGCLKBUF),.T3I3(NET_10),.TB3S(GND),.C3Z(NET_594),.Q3Z(tcdm_result_p1[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_O16_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B0I0(tcdm_rdata_p1_int[19]),.B0I1(tcdm_rdata_p3_int[19]),.B0I2(NET_110),.B0I3(NET_125),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[17]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p1_int[19]),.T0I1(tcdm_rdata_p3_int[19]),.T0I2(NET_110),.T0I3(NET_125),.TB0S(NET_10),.C0Z(NET_382),.Q0Z(tcdm_result_p3[17]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B1I0(tcdm_result_p3[19]),.B1I1(NET_96),.B1I2(fpgaio_out_dup_0[51]),.B1I3(NET_99),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[51]),.T1I1(NET_99),.T1I2(tcdm_result_p3[19]),.T1I3(NET_96),.TB1S(NET_376),.C1Z(NET_373),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_O16_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_125),.B2I1(tcdm_rdata_p3_int[17]),.B2I2(NET_110),.B2I3(tcdm_rdata_p1_int[17]),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[19]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_125),.T2I1(tcdm_rdata_p3_int[17]),.T2I2(NET_110),.T2I3(tcdm_rdata_p1_int[17]),.TB2S(NET_10),.C2Z(NET_345),.Q2Z(tcdm_result_p3[19]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O16_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.B3I0(lint_ADDR_int[3]),.B3I1(lint_ADDR_int[5]),.B3I2(lint_ADDR_int[4]),.B3I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[4]),.T3I1(lint_ADDR_int[11]),.T3I2(lint_ADDR_int[3]),.T3I3(lint_ADDR_int[5]),.TB3S(lint_ADDR_int[6]),.C3Z(NET_125),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_O17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O17_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B1I0(NET_125),.B1I1(NET_110),.B1I2(tcdm_rdata_p3_int[29]),.B1I3(tcdm_rdata_p1_int[29]),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[26]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p3_int[29]),.T1I1(tcdm_rdata_p1_int[29]),.T1I2(NET_125),.T1I3(NET_110),.TB1S(NET_10),.C1Z(NET_581),.Q1Z(tcdm_result_p3[26]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_O17_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_125),.B2I1(NET_110),.B2I2(tcdm_rdata_p1_int[28]),.B2I3(tcdm_rdata_p3_int[28]),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_125),.T2I1(NET_110),.T2I2(tcdm_rdata_p1_int[28]),.T2I3(tcdm_rdata_p3_int[28]),.TB2S(NET_10),.C2Z(NET_563),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_O17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(tcdm_result_p3[26]),.B3I1(NET_96),.B3I2(NET_99),.B3I3(fpgaio_out_dup_0[58]),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[29]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_99),.T3I1(fpgaio_out_dup_0[58]),.T3I2(tcdm_result_p3[26]),.T3I3(NET_96),.TB3S(NET_522),.C3Z(NET_519),.Q3Z(tcdm_result_p3[29]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_O18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(tcdm_result_p3[28]),.B0I1(NET_96),.B0I2(fpgaio_out_dup_0[60]),.B0I3(NET_99),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[28]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p3[28]),.T0I1(NET_96),.T0I2(fpgaio_out_dup_0[60]),.T0I3(NET_99),.TB0S(NET_557),.C0Z(NET_554),.Q0Z(tcdm_result_p3[28]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B1I0(tcdm_result_p3[22]),.B1I1(NET_99),.B1I2(fpgaio_out_dup_0[54]),.B1I3(NET_96),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[54]),.T1I1(NET_96),.T1I2(tcdm_result_p3[22]),.T1I3(NET_99),.TB1S(NET_430),.C1Z(NET_427),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_O18_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B2I0(tcdm_rdata_p1_int[21]),.B2I1(NET_125),.B2I2(NET_110),.B2I3(tcdm_rdata_p3_int[21]),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[21]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p1_int[21]),.T2I1(NET_125),.T2I2(NET_110),.T2I3(tcdm_rdata_p3_int[21]),.TB2S(NET_10),.C2Z(NET_418),.Q2Z(tcdm_result_p3[21]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B3I0(tcdm_result_p3[21]),.B3I1(fpgaio_out_dup_0[53]),.B3I2(NET_99),.B3I3(NET_96),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_99),.T3I1(NET_96),.T3I2(tcdm_result_p3[21]),.T3I3(fpgaio_out_dup_0[53]),.TB3S(NET_412),.C3Z(NET_409),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_O19_0 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(GND),.B0I1(lint_ADDR_int[11]),.B0I2(GND),.B0I3(lint_ADDR_int[6]),.T0I0(GND),.T0I1(NET_69),.T0I2(NET_75),.T0I3(NET_77),.TB0S(GND),.B0Z(NET_77),.C0Z(NET_66),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_O19_1 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(GND),.T1I1(lint_ADDR_int[11]),.T1I2(NET_75),.T1I3(lint_ADDR_int[2]),.C1Z(NET_76),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O19_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000001),.B2I0(GND),.B2I1(lint_ADDR_int[5]),.B2I2(GND),.B2I3(lint_ADDR_int[7]),.T2I0(lint_ADDR_int[4]),.T2I1(lint_ADDR_int[13]),.T2I2(GND),.T2I3(lint_ADDR_int[10]),.TB2S(GND),.B2Z(NET_75),.C2Z(NET_150),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_O19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_75),.B3I1(NET_77),.B3I2(NET_149),.B3I3(NET_71),.T3I0(NET_149),.T3I1(NET_71),.T3I2(NET_75),.T3I3(NET_77),.TB3S(NET_150),.C3Z(NET_147),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_O20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O20_1 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(GND),.T1I1(lint_ADDR_int[2]),.T1I2(lint_ADDR_int[3]),.T1I3(GND),.C1Z(NET_134),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O23_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_141),.T1I1(NET_142),.T1I2(NET_646),.T1I3(GND),.TB1S(GND),.C1Z(nx53672z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_O23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O23_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_141),.T3I1(NET_142),.T3I2(NET_140),.T3I3(GND),.C3Z(nx14650z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O27_3 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int[13]),.T3I1(NET_252),.T3I2(NET_65),.T3I3(NET_143),.TB3S(GND),.C3Z(nx30664z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_O28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[6]),.Q2EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_waddr_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O32_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[3]),.Q0EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_rdata_int[11]),.T0I1(NET_44_CAND4_BLSBR_15_tpGCLKBUF),.T0I2(m1_coef_rdata_int[11]),.T0I3(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.TB0S(GND),.C0Z(NET_203),.Q0Z(m1_coef_waddr_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O32_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(m1_oper1_rdata_int[14]),.T1I1(NET_44_CAND4_BLSBR_15_tpGCLKBUF),.T1I2(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.T1I3(m1_coef_rdata_int[14]),.C1Z(NET_263),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O32_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_oper1_rdata_int[5]),.B2I1(NET_44_CAND4_BLSBR_15_tpGCLKBUF),.B2I2(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.B2I3(m1_coef_rdata_int[5]),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_44_CAND4_BLSBR_15_tpGCLKBUF),.T2I1(m1_coef_rdata_int[10]),.T2I2(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.T2I3(m1_oper1_rdata_int[10]),.TB2S(GND),.B2Z(NET_657),.C2Z(NET_184),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_O32_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(m1_oper1_rdata_int[15]),.T3I1(m1_coef_rdata_int[15]),.T3I2(NET_44_CAND4_BLSBR_15_tpGCLKBUF),.T3I3(NET_43_CAND3_BLSBR_15_tpGCLKBUF),.TB3S(GND),.C3Z(NET_302),.Q3Z(m1_coef_wdata_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_P1_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[5]),.Q0EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.T0I0(NET_41),.T0I1(m0_coef_rdata_int[18]),.T0I2(NET_46_CAND1_TLSTR_16_tpGCLKBUF),.T0I3(m0_oper1_rdata_int[18]),.TB0S(GND),.C0Z(NET_366),.Q0Z(m0_coef_waddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[4]),.Q1EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_waddr_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[10]),.Q2EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_waddr_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P1_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.T3I0(NET_46_CAND1_TLSTR_16_tpGCLKBUF),.T3I1(NET_41),.T3I2(m0_oper1_rdata_int[29]),.T3I3(m0_coef_rdata_int[29]),.C3Z(NET_584),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[8]),.Q0EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_waddr_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[1]),.Q1EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_waddr_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[3]),.Q2EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_waddr_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[11]),.Q3EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_waddr_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[2]),.Q0EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_waddr_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[9]),.Q1EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_waddr_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[7]),.Q2EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_waddr_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(NET_762),.Q3EN(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_we_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_outsel_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_reset_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_outsel_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_outsel_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P9_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[3]),.T1I1(lint_ADDR_int[4]),.T1I2(lint_ADDR_int[5]),.T1I3(lint_ADDR_int[6]),.C1Z(NET_15),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_P9_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND),.C2Z(NET_762),.Q2Z(m0_m1_rnd_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_P9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P11_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[17]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(m0_m1_rnd_dup_0),.T0I1(NET_51),.T0I2(NET_63),.T0I3(tcdm_result_p3[16]),.TB0S(GND),.C0Z(NET_324),.Q0Z(m0_m1_clr_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P11_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T1I0(NET_51),.T1I1(NET_63),.T1I2(m0_m1_reset_dup_0),.T1I3(tcdm_result_p3[31]),.TB1S(GND),.C1Z(NET_614),.Q1Z(m0_m1_control[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_P11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P11_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T3I0(NET_51),.T3I1(NET_63),.T3I2(tcdm_result_p3[20]),.T3I3(m0_m1_control[20]),.TB3S(GND),.C3Z(NET_398),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_P12_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[31]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p0[25]),.T0I1(NET_34),.T0I2(NET_13),.T0I3(tcdm_rdata_p3_int[25]),.TB0S(GND),.C0Z(NET_512),.Q0Z(tcdm_result_p3[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[16]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p3[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_34),.B2I1(tcdm_rdata_p3_int[20]),.B2I2(NET_13),.B2I3(tcdm_result_p0[20]),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[25]),.Q2EN(tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.B2Z(NET_402),.Q2Z(tcdm_result_p0[25]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[20]),.Q3EN(tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P13_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_34),.B0I1(NET_13),.B0I2(tcdm_rdata_p3_int[30]),.B0I3(tcdm_result_p0[30]),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[27]),.Q0EN(tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(NET_34),.T0I1(tcdm_rdata_p3_int[31]),.T0I2(NET_13),.T0I3(tcdm_result_p0[31]),.TB0S(GND),.B0Z(NET_600),.C0Z(NET_618),.Q0Z(tcdm_result_p0[27]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P13_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[30]),.Q1EN(tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p3_int[27]),.T1I1(tcdm_result_p0[27]),.T1I2(NET_13),.T1I3(NET_34),.TB1S(GND),.C1Z(NET_547),.Q1Z(tcdm_result_p0[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_P13_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000001000000000),.B2I0(NET_14),.B2I1(GND),.B2I2(GND),.B2I3(NET_15_CAND5_TLSBR_16_tpGCLKBUF),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[16]),.Q2EN(tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T2I0(NET_7),.T2I1(GND),.T2I2(GND),.T2I3(NET_49),.TB2S(GND),.B2Z(NET_13),.C2Z(NET_51),.Q2Z(tcdm_result_p0[16]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_P13_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[31]),.Q3EN(tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p0[16]),.T3I1(tcdm_rdata_p3_int[16]),.T3I2(NET_13),.T3I3(NET_34),.C3Z(NET_328),.Q3Z(tcdm_result_p0[31]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000010000),.B0I0(lint_ADDR_int[8]),.B0I1(apb_fsm[0]),.B0I2(lint_ADDR_int[7]),.B0I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[8]),.T0I1(apb_fsm[0]),.T0I2(lint_ADDR_int[7]),.T0I3(lint_ADDR_int[11]),.TB0S(lint_ADDR_int[2]),.C0Z(NET_101),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P14_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B1I0(tcdm_result_p1[24]),.B1I1(NET_101),.B1I2(tcdm_result_p0[24]),.B1I3(NET_89),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[24]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p0[24]),.T1I1(NET_89),.T1I2(tcdm_result_p1[24]),.T1I3(NET_101),.TB1S(NET_15_CAND5_TLSBR_16_tpGCLKBUF),.C1Z(NET_487),.Q1Z(tcdm_result_p1[24]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_P14_2 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[24]),.Q2EN(tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[8]),.T2I1(apb_fsm[0]),.T2I2(lint_ADDR_int[7]),.T2I3(lint_ADDR_int[2]),.TB2S(GND),.C2Z(NET_49),.Q2Z(tcdm_result_p0[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_P14_3 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[8]),.T3I1(apb_fsm[0]),.T3I2(lint_ADDR_int[2]),.T3I3(lint_ADDR_int[7]),.C3Z(NET_14),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P15_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(tcdm_result_p1[18]),.B0I1(tcdm_result_p0[18]),.B0I2(NET_101),.B0I3(NET_89),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[18]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p1[18]),.T0I1(tcdm_result_p0[18]),.T0I2(NET_101),.T0I3(NET_89),.TB0S(NET_15_CAND5_TLSBR_16_tpGCLKBUF),.C0Z(NET_357),.Q0Z(tcdm_result_p1[18]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[22]),.Q1EN(tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000100000000),.B2I0(GND),.B2I1(apb_fsm[0]),.B2I2(lint_ADDR_int[11]),.B2I3(lint_ADDR_int[8]),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[18]),.Q2EN(tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.B2Z(NET_87),.Q2Z(tcdm_result_p0[18]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P15_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B3I0(tcdm_result_p0[22]),.B3I1(tcdm_result_p1[22]),.B3I2(NET_89),.B3I3(NET_101),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[22]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T3I0(NET_89),.T3I1(NET_101),.T3I2(tcdm_result_p0[22]),.T3I3(tcdm_result_p1[22]),.TB3S(NET_15_CAND5_TLSBR_16_tpGCLKBUF),.C3Z(NET_430),.Q3Z(tcdm_result_p1[22]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_P16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001000000000000),.B0I0(GND),.B0I1(GND),.B0I2(NET_101),.B0I3(NET_7),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.B0Z(NET_99),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P16_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(tcdm_rdata_p3_int[18]),.B1I1(NET_125),.B1I2(NET_110),.B1I3(tcdm_rdata_p1_int[18]),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T1I0(NET_110),.T1I1(tcdm_rdata_p1_int[18]),.T1I2(tcdm_rdata_p3_int[18]),.T1I3(NET_125),.TB1S(NET_10),.C1Z(NET_363),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_P16_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_125),.B2I1(tcdm_rdata_p3_int[7]),.B2I2(NET_110),.B2I3(tcdm_rdata_p1_int[7]),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T2I0(NET_125),.T2I1(tcdm_rdata_p3_int[7]),.T2I2(NET_110),.T2I3(tcdm_rdata_p1_int[7]),.TB2S(NET_10),.C2Z(NET_478),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_P16_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B3I0(NET_110),.B3I1(NET_125),.B3I2(tcdm_rdata_p1_int[6]),.B3I3(tcdm_rdata_p3_int[6]),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[18]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p1_int[6]),.T3I1(tcdm_rdata_p3_int[6]),.T3I2(NET_110),.T3I3(NET_125),.TB3S(NET_10),.C3Z(NET_644),.Q3Z(tcdm_result_p3[18]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_P18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P18_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B1I0(NET_110),.B1I1(tcdm_rdata_p1_int[24]),.B1I2(NET_125),.B1I3(tcdm_rdata_p3_int[24]),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T1I0(NET_125),.T1I1(tcdm_rdata_p3_int[24]),.T1I2(NET_110),.T1I3(tcdm_rdata_p1_int[24]),.TB1S(NET_10),.C1Z(NET_493),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_P18_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B2I0(tcdm_rdata_p1_int[22]),.B2I1(tcdm_rdata_p3_int[22]),.B2I2(NET_125),.B2I3(NET_110),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[24]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p1_int[22]),.T2I1(tcdm_rdata_p3_int[22]),.T2I2(NET_125),.T2I3(NET_110),.TB2S(NET_10),.C2Z(NET_436),.Q2Z(tcdm_result_p3[24]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_P18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[22]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p3[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000100000000),.B0I0(GND),.B0I1(apb_fsm[0]),.B0I2(GND),.B0I3(lint_ADDR_int[8]),.B0Z(NET_19),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P19_1 (.tFragBitInfo(16'b0011011100111111),.bFragBitInfo(16'b0000000011111111),.B1I0(NET_76),.B1I1(NET_172),.B1I2(NET_77),.B1I3(NET_69),.T1I0(NET_77),.T1I1(NET_69),.T1I2(NET_76),.T1I3(NET_172),.TB1S(NET_148),.C1Z(NET_620),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_P19_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000001000),.B2I0(NET_77),.B2I1(NET_69),.B2I2(GND),.B2I3(GND),.T2I0(NET_65),.T2I1(GND),.T2I2(GND),.T2I3(NET_148),.TB2S(GND),.B2Z(NET_132),.C2Z(NET_173),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_P19_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_76),.T3I1(NET_69),.T3I2(GND),.T3I3(GND),.C3Z(NET_68),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[2]),.Q0EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_waddr_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(NET_762),.Q2EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_we_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[9]),.Q3EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_waddr_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[0]),.Q0EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_waddr_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[5]),.Q1EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_waddr_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[11]),.Q2EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_waddr_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[4]),.Q3EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_waddr_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[7]),.Q0EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_waddr_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[8]),.Q1EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_waddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[1]),.Q2EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_waddr_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_16_padClk),.QRT(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_waddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_46),.B0I1(m0_oper1_rdata_int[16]),.B0I2(NET_41),.B0I3(m0_coef_rdata_int[16]),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.B0Z(NET_325),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[4]),.Q1EN(nx32231z1_CAND2_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_raddr_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q1_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_46),.B2I1(m0_coef_rdata_int[20]),.B2I2(m0_oper1_rdata_int[20]),.B2I3(NET_41),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.T2I0(NET_46),.T2I1(m0_oper1_rdata_int[25]),.T2I2(NET_41),.T2I3(m0_coef_rdata_int[25]),.TB2S(GND),.B2Z(NET_399),.C2Z(NET_509),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_Q1_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[6]),.Q3EN(nx32231z1_CAND2_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.T3I0(NET_46),.T3I1(NET_41),.T3I2(m0_oper1_rdata_int[19]),.T3I3(m0_coef_rdata_int[19]),.TB3S(GND),.C3Z(NET_385),.Q3Z(m0_coef_raddr_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Q2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[9]),.Q0EN(nx32231z1_CAND2_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_raddr_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[7]),.Q1EN(nx32231z1_CAND2_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_raddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[8]),.Q2EN(nx32231z1_CAND2_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_raddr_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[11]),.Q3EN(nx32231z1_CAND2_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_raddr_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[20]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p3[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q13_0 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T0I0(NET_49_CAND4_TRSBL_17_tpGCLKBUF),.T0I1(NET_15),.T0I2(GND),.T0I3(GND),.TB0S(GND),.C0Z(NET_50),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q13_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[27]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[2]),.T3I1(NET_15),.T3I2(NET_19),.T3I3(lint_ADDR_int[7]),.TB3S(GND),.C3Z(NET_52),.Q3Z(tcdm_result_p3[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Q14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001000),.B0I0(NET_15),.B0I1(NET_10),.B0I2(GND),.B0I3(GND),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B0Z(NET_35),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q14_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B1I0(tcdm_result_p1[23]),.B1I1(NET_89),.B1I2(NET_101),.B1I3(tcdm_result_p0[23]),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[23]),.Q1EN(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T1I0(NET_101),.T1I1(tcdm_result_p0[23]),.T1I2(tcdm_result_p1[23]),.T1I3(NET_89),.TB1S(NET_15),.C1Z(NET_448),.Q1Z(tcdm_result_p1[23]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_Q14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[23]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p0[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q14_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T3I0(NET_7_CAND3_TRSBL_17_tpGCLKBUF),.T3I1(NET_10),.T3I2(GND),.T3I3(GND),.C3Z(NET_34),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_Q15_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(tcdm_result_p1[28]),.B0I1(NET_89),.B0I2(NET_101),.B0I3(tcdm_result_p0[28]),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[28]),.Q0EN(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p1[28]),.T0I1(NET_89),.T0I2(NET_101),.T0I3(tcdm_result_p0[28]),.TB0S(NET_15),.C0Z(NET_557),.Q0Z(tcdm_result_p1[28]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q15_1 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[28]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T1I0(NET_7_CAND3_TRSBL_17_tpGCLKBUF),.T1I1(NET_89),.T1I2(GND),.T1I3(GND),.TB1S(GND),.C1Z(NET_82),.Q1Z(tcdm_result_p0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_Q15_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B2I0(tcdm_result_p0[26]),.B2I1(NET_89),.B2I2(NET_101),.B2I3(tcdm_result_p1[26]),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[26]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p0[26]),.T2I1(NET_89),.T2I2(NET_101),.T2I3(tcdm_result_p1[26]),.TB2S(NET_15),.C2Z(NET_522),.Q2Z(tcdm_result_p0[26]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_Q15_3 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[26]),.Q3EN(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_101),.T3I2(GND),.T3I3(NET_15),.C3Z(NET_100),.Q3Z(tcdm_result_p1[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_Q17_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_100),.B0I1(tcdm_result_p1[0]),.B0I2(NET_99),.B0I3(tcdm_result_p3[0]),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[0]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND1_BRSTL_17_tpGCLKBUF),.QST(GND),.T0I0(NET_100),.T0I1(NET_99),.T0I2(tcdm_result_p1[12]),.T0I3(tcdm_result_p3[12]),.TB0S(GND),.B0Z(NET_91),.C0Z(NET_218),.Q0Z(tcdm_result_p1[0]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q17_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B1I0(tcdm_rdata_p3_int[12]),.B1I1(NET_125_CAND3_BRSTL_17_tpGCLKBUF),.B1I2(tcdm_rdata_p1_int[12]),.B1I3(NET_110_CAND4_BRSTL_17_tpGCLKBUF),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[0]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND1_BRSTL_17_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p1_int[12]),.T1I1(NET_110_CAND4_BRSTL_17_tpGCLKBUF),.T1I2(tcdm_rdata_p3_int[12]),.T1I3(NET_125_CAND3_BRSTL_17_tpGCLKBUF),.TB1S(NET_10),.C1Z(NET_232),.Q1Z(tcdm_result_p3[0]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_Q17_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B2I0(tcdm_rdata_p3_int[0]),.B2I1(NET_110_CAND4_BRSTL_17_tpGCLKBUF),.B2I2(NET_125_CAND3_BRSTL_17_tpGCLKBUF),.B2I3(tcdm_rdata_p1_int[0]),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[12]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND1_BRSTL_17_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p3_int[0]),.T2I1(NET_110_CAND4_BRSTL_17_tpGCLKBUF),.T2I2(NET_125_CAND3_BRSTL_17_tpGCLKBUF),.T2I3(tcdm_rdata_p1_int[0]),.TB2S(NET_10),.C2Z(NET_130),.Q2Z(tcdm_result_p1[12]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_Q17_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001010100111111),.B3I0(NET_125_CAND3_BRSTL_17_tpGCLKBUF),.B3I1(tcdm_rdata_p3_int[2]),.B3I2(NET_110_CAND4_BRSTL_17_tpGCLKBUF),.B3I3(tcdm_rdata_p1_int[2]),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[12]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND1_BRSTL_17_tpGCLKBUF),.QST(GND),.T3I0(NET_110_CAND4_BRSTL_17_tpGCLKBUF),.T3I1(tcdm_rdata_p1_int[2]),.T3I2(NET_125_CAND3_BRSTL_17_tpGCLKBUF),.T3I3(tcdm_rdata_p3_int[2]),.TB3S(NET_10),.C3Z(NET_725),.Q3Z(tcdm_result_p3[12]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Q18_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001001101011111),.B0I0(tcdm_rdata_p3_int[23]),.B0I1(NET_125_CAND3_BRSTL_17_tpGCLKBUF),.B0I2(NET_110_CAND4_BRSTL_17_tpGCLKBUF),.B0I3(tcdm_rdata_p1_int[23]),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND1_BRSTL_17_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p3_int[23]),.T0I1(NET_125_CAND3_BRSTL_17_tpGCLKBUF),.T0I2(NET_110_CAND4_BRSTL_17_tpGCLKBUF),.T0I3(tcdm_rdata_p1_int[23]),.TB0S(NET_10),.C0Z(NET_454),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND1_BRSTL_17_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND1_BRSTL_17_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q18_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0000011101110111),.B3I0(tcdm_rdata_p1_int[26]),.B3I1(NET_125_CAND3_BRSTL_17_tpGCLKBUF),.B3I2(tcdm_rdata_p3_int[26]),.B3I3(NET_110_CAND4_BRSTL_17_tpGCLKBUF),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[23]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND1_BRSTL_17_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p3_int[26]),.T3I1(NET_110_CAND4_BRSTL_17_tpGCLKBUF),.T3I2(tcdm_rdata_p1_int[26]),.T3I3(NET_125_CAND3_BRSTL_17_tpGCLKBUF),.TB3S(NET_10),.C3Z(NET_528),.Q3Z(tcdm_result_p3[23]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Q31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[11]),.Q0EN(nx14650z1_CAND2_BRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND1_BRSBL_17_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_raddr_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[4]),.Q1EN(nx14650z1_CAND2_BRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND1_BRSBL_17_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[6]),.Q2EN(nx14650z1_CAND2_BRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND1_BRSBL_17_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_raddr_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[5]),.Q3EN(nx14650z1_CAND2_BRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND1_BRSBL_17_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_raddr_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[7]),.Q0EN(nx14650z1_CAND2_BRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND1_BRSBL_17_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_raddr_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[10]),.Q1EN(nx14650z1_CAND2_BRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND1_BRSBL_17_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[9]),.Q2EN(nx14650z1_CAND2_BRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND1_BRSBL_17_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_raddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[8]),.Q3EN(nx14650z1_CAND2_BRSBL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND1_BRSBL_17_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_raddr_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[1]),.Q0EN(nx32231z1_CAND2_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_raddr_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[5]),.Q1EN(nx32231z1_CAND2_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_raddr_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[0]),.Q2EN(nx32231z1_CAND2_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_raddr_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx32231z1_CAND2_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_raddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[3]),.Q0EN(nx32231z1_CAND2_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_raddr_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[2]),.Q3EN(nx32231z1_CAND2_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_raddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100000000000),.B1I0(NET_139),.B1I1(lint_ADDR_int[2]),.B1I2(lint_ADDR_int[3]),.B1I3(NET_132),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[3]),.T1I1(NET_132),.T1I2(NET_139),.T1I3(lint_ADDR_int[2]),.TB1S(lint_ADDR_int[4]),.Q1Z(m0_m1_clken_dup_0),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_R8_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T2I0(NET_138),.T2I1(NET_132),.T2I2(lint_ADDR_int[4]),.T2I3(NET_139),.TB2S(GND),.Q2Z(m0_m0_clken_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_R8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B2I0(lint_ADDR_int[5]),.B2I1(lint_ADDR_int[7]),.B2I2(GND),.B2I3(NET_65),.B2Z(NET_139),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R12_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_48),.B2I1(m0_m1_dataout_int[20]),.B2I2(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.B2I3(tcdm_result_p2[20]),.T2I0(m0_m1_dataout_int[25]),.T2I1(tcdm_result_p2[25]),.T2I2(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.T2I3(NET_48),.TB2S(GND),.B2Z(NET_387),.C2Z(NET_497),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_R12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R13_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B0I0(m0_m1_dataout_int[16]),.B0I1(tcdm_result_p2[16]),.B0I2(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.B0I3(NET_48),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[16]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(m0_m1_dataout_int[30]),.T0I1(tcdm_result_p2[30]),.T0I2(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.T0I3(NET_48),.TB0S(GND),.B0Z(NET_312),.C0Z(NET_585),.Q0Z(tcdm_result_p2[16]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R13_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[25]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p2[31]),.T1I1(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.T1I2(m0_m1_dataout_int[31]),.T1I3(NET_48),.TB1S(GND),.C1Z(NET_603),.Q1Z(tcdm_result_p2[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_R13_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[31]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p2[27]),.T2I1(m0_m1_dataout_int[27]),.T2I2(NET_52_CAND2_TRSBL_18_tpGCLKBUF),.T2I3(NET_48),.TB2S(GND),.C2Z(NET_532),.Q2Z(tcdm_result_p2[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_R13_3 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[20]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_14),.T3I2(NET_7_CAND3_TRSBL_18_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.C3Z(NET_48),.Q3Z(tcdm_result_p2[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_R14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[27]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p2[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[30]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R15_0 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0000000000000000),.T0I0(lint_ADDR_int[7]),.T0I1(NET_87),.T0I2(lint_ADDR_int[2]),.T0I3(NET_15),.TB0S(GND),.C0Z(NET_86),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_R15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[6]),.Q0EN(tcdm_valid_p1_int_CAND5_TRSBL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p1[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R16_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[7]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[2]),.T1I1(lint_ADDR_int[7]),.T1I2(NET_87),.T1I3(NET_7_CAND3_TRSBL_18_tpGCLKBUF),.C1Z(NET_83),.Q1Z(tcdm_result_p3[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_R16_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[6]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(NET_99),.T2I1(NET_100),.T2I2(tcdm_result_p1[7]),.T2I3(tcdm_result_p3[7]),.TB2S(GND),.C2Z(NET_464),.Q2Z(tcdm_result_p3[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_R16_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[7]),.Q3EN(tcdm_valid_p1_int_CAND5_TRSBL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T3I0(NET_99),.T3I1(tcdm_result_p1[6]),.T3I2(tcdm_result_p3[6]),.T3I3(NET_100),.C3Z(NET_630),.Q3Z(tcdm_result_p1[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_R17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_99),.B0I1(tcdm_result_p1[2]),.B0I2(tcdm_result_p3[2]),.B0I3(NET_100),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[2]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND1_BRSTL_18_tpGCLKBUF),.QST(GND),.B0Z(NET_711),.Q0Z(tcdm_result_p1[2]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R17_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND1_BRSTL_18_tpGCLKBUF),.QST(GND),.T1I0(NET_83_CAND2_BRSTL_18_tpGCLKBUF),.T1I1(m1_m1_dataout_int[29]),.T1I2(NET_86),.T1I3(m0_m1_dataout_int[29]),.C1Z(NET_571),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_R17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[2]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND1_BRSTL_18_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R17_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND1_BRSTL_18_tpGCLKBUF),.QST(GND),.T3I0(NET_83_CAND2_BRSTL_18_tpGCLKBUF),.T3I1(m1_m1_dataout_int[26]),.T3I2(NET_86),.T3I3(m0_m1_dataout_int[26]),.C3Z(NET_518),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_R18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R18_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_m1_dataout_int[28]),.T1I1(NET_83_CAND2_BRSTL_18_tpGCLKBUF),.T1I2(m1_m1_dataout_int[28]),.T1I3(NET_86),.TB1S(GND),.C1Z(NET_553),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_R18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_m1_dataout_int[24]),.B2I1(NET_83_CAND2_BRSTL_18_tpGCLKBUF),.B2I2(m0_m1_dataout_int[24]),.B2I3(NET_86),.B2Z(NET_483),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND1_BRSTL_18_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND1_BRSTL_18_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000010000000),.B2I0(NET_139),.B2I1(NET_132),.B2I2(lint_ADDR_int[3]),.B2I3(lint_ADDR_int[2]),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND1_BRSTL_18_tpGCLKBUF),.QST(GND),.T2I0(NET_139),.T2I1(NET_132),.T2I2(lint_ADDR_int[3]),.T2I3(lint_ADDR_int[2]),.TB2S(lint_ADDR_int[4]),.Q2Z(m1_m0_clken_dup_0),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_R20_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND1_BRSTL_18_tpGCLKBUF),.QST(GND),.T3I0(NET_139),.T3I1(NET_132),.T3I2(NET_134),.T3I3(lint_ADDR_int[4]),.TB3S(GND),.Q3Z(m1_m1_clken_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_R31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND1_BRSBL_18_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND1_BRSBL_18_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND1_BRSBL_18_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[2]),.Q3EN(nx14650z1_CAND2_BRSBL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND1_BRSBL_18_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_raddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[1]),.Q0EN(nx14650z1_CAND2_BRSBL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND1_BRSBL_18_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_raddr_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[0]),.Q1EN(nx14650z1_CAND2_BRSBL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND1_BRSBL_18_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND1_BRSBL_18_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[3]),.Q3EN(nx14650z1_CAND2_BRSBL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND1_BRSBL_18_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_raddr_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[5]),.Q0EN(tcdm_valid_p1_int_CAND5_TRSBL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p1[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S12_2 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0000000000101010),.B2I0(NET_756),.B2I1(m0_m1_dataout_int[5]),.B2I2(NET_52_CAND2_TRSBL_19_tpGCLKBUF),.B2I3(tcdm_result_p1[5]),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T2I0(NET_756),.T2I1(m0_m1_dataout_int[5]),.T2I2(NET_52_CAND2_TRSBL_19_tpGCLKBUF),.T2I3(tcdm_result_p1[5]),.TB2S(NET_50),.C2Z(NET_757),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_S12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S13_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[5]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T0I0(NET_34),.T0I1(tcdm_rdata_p3_int[5]),.T0I2(tcdm_rdata_p1_int[5]),.T0I3(NET_35),.TB0S(GND),.C0Z(NET_653),.Q0Z(tcdm_result_p3[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S13_2 (.tFragBitInfo(16'b0101111111111111),.bFragBitInfo(16'b0001111100111111),.B2I0(tcdm_result_p3[5]),.B2I1(tcdm_result_p2[5]),.B2I2(NET_7_CAND3_TRSBL_19_tpGCLKBUF),.B2I3(NET_49_CAND4_TRSBL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p3[5]),.T2I1(tcdm_result_p2[5]),.T2I2(NET_7_CAND3_TRSBL_19_tpGCLKBUF),.T2I3(NET_49_CAND4_TRSBL_19_tpGCLKBUF),.TB2S(NET_14),.C2Z(NET_756),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_S13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S14_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_146),.T2I1(lint_ADDR_int[5]),.T2I2(lint_ADDR_int[6]),.T2I3(NET_145),.TB2S(GND),.C2Z(nx49871z1),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S15_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T1I0(NET_85),.T1I1(m1_ram_control[2]),.T1I2(m0_m1_dataout_int[2]),.T1I3(NET_86),.TB1S(GND),.C1Z(NET_709),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_S15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.Q2Z(m1_ram_control[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_S15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S16_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_83),.T1I1(m0_m1_dataout_int[19]),.T1I2(m1_m1_dataout_int[19]),.T1I3(NET_86),.C1Z(NET_372),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_83),.B2I1(m0_m1_dataout_int[18]),.B2I2(NET_86),.B2I3(m1_m1_dataout_int[18]),.B2Z(NET_353),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_S16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[5]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p2[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[2]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S17_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(m0_m1_dataout_int[22]),.T2I1(NET_83_CAND2_BRSTL_19_tpGCLKBUF),.T2I2(NET_86),.T2I3(m1_m1_dataout_int[22]),.TB2S(GND),.C2Z(NET_426),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_S17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B3I0(tcdm_result_p2[2]),.B3I1(NET_82),.B3I2(m1_m1_dataout_int[2]),.B3I3(NET_83_CAND2_BRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF),.QST(GND),.T3I0(m1_m1_dataout_int[2]),.T3I1(NET_83_CAND2_BRSTL_19_tpGCLKBUF),.T3I2(tcdm_result_p2[2]),.T3I3(NET_82),.TB3S(NET_709),.C3Z(NET_707),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_S18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S18_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_m1_dataout_int[23]),.T1I1(m1_m1_dataout_int[23]),.T1I2(NET_86),.T1I3(NET_83_CAND2_BRSTL_19_tpGCLKBUF),.C1Z(NET_444),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_m1_dataout_int[21]),.B2I1(NET_83_CAND2_BRSTL_19_tpGCLKBUF),.B2I2(NET_86),.B2I3(m0_m1_dataout_int[21]),.B2Z(NET_408),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_S18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_T12_0 (.tFragBitInfo(16'b0111000001110000),.bFragBitInfo(16'b0000000001110000),.B0I0(m0_m1_dataout_int[14]),.B0I1(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.B0I2(NET_737),.B0I3(tcdm_result_p1[14]),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T0I0(m0_m1_dataout_int[14]),.T0I1(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.T0I2(NET_737),.T0I3(tcdm_result_p1[14]),.TB0S(NET_50),.C0Z(NET_738),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T12_1 (.tFragBitInfo(16'b0011111100000000),.bFragBitInfo(16'b0000010000001100),.B1I0(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.B1I1(NET_733),.B1I2(tcdm_result_p1[11]),.B1I3(m0_m1_dataout_int[11]),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[14]),.Q1EN(tcdm_valid_p1_int_CAND5_TRSBL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p1[11]),.T1I1(m0_m1_dataout_int[11]),.T1I2(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.T1I3(NET_733),.TB1S(NET_50),.C1Z(NET_734),.Q1Z(tcdm_result_p1[14]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_T12_2 (.tFragBitInfo(16'b0111000001110000),.bFragBitInfo(16'b0000000001110000),.B2I0(m0_m1_dataout_int[15]),.B2I1(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.B2I2(NET_741),.B2I3(tcdm_result_p1[15]),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T2I0(m0_m1_dataout_int[15]),.T2I1(NET_52_CAND2_TRSBL_20_tpGCLKBUF),.T2I2(NET_741),.T2I3(tcdm_result_p1[15]),.TB2S(NET_50),.C2Z(NET_742),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_T12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[15]),.Q3EN(tcdm_valid_p1_int_CAND5_TRSBL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p1[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_T14_0 (.tFragBitInfo(16'b0111111101111111),.bFragBitInfo(16'b0000111101111111),.B0I0(tcdm_result_p3[14]),.B0I1(NET_49_CAND4_TRSBL_20_tpGCLKBUF),.B0I2(NET_7_CAND3_TRSBL_20_tpGCLKBUF),.B0I3(tcdm_result_p2[14]),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[14]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p3[14]),.T0I1(NET_49_CAND4_TRSBL_20_tpGCLKBUF),.T0I2(NET_7_CAND3_TRSBL_20_tpGCLKBUF),.T0I3(tcdm_result_p2[14]),.TB0S(NET_14),.C0Z(NET_737),.Q0Z(tcdm_result_p3[14]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T14_1 (.tFragBitInfo(16'b0111011111111111),.bFragBitInfo(16'b0011011101110111),.B1I0(tcdm_result_p2[15]),.B1I1(NET_7_CAND3_TRSBL_20_tpGCLKBUF),.B1I2(tcdm_result_p3[15]),.B1I3(NET_49_CAND4_TRSBL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p3[15]),.T1I1(NET_49_CAND4_TRSBL_20_tpGCLKBUF),.T1I2(tcdm_result_p2[15]),.T1I3(NET_7_CAND3_TRSBL_20_tpGCLKBUF),.TB1S(NET_14),.C1Z(NET_741),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_T14_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[15]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p1_int[15]),.T2I1(tcdm_rdata_p3_int[15]),.T2I2(NET_35),.T2I3(NET_34),.TB2S(GND),.C2Z(NET_298),.Q2Z(tcdm_result_p3[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_T14_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p3_int[14]),.T3I1(NET_34),.T3I2(NET_35),.T3I3(tcdm_rdata_p1_int[14]),.C3Z(NET_259),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_T15_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T0I0(m0_m1_dataout_int[12]),.T0I1(NET_85),.T0I2(NET_86),.T0I3(m1_ram_control[12]),.TB0S(GND),.C0Z(NET_216),.Q0Z(m1_ram_control[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.Q1Z(m1_ram_control[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T15_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B2I0(m0_m1_dataout_int[7]),.B2I1(m1_ram_control[7]),.B2I2(NET_86),.B2I3(NET_85),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T2I0(m1_ram_control[0]),.T2I1(m0_m1_dataout_int[0]),.T2I2(NET_86),.T2I3(NET_85),.TB2S(GND),.B2Z(NET_462),.C2Z(NET_84),.Q2Z(m1_ram_control[0]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_T15_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T3I0(m0_m1_dataout_int[6]),.T3I1(NET_85),.T3I2(NET_86),.T3I3(m1_ram_control[6]),.C3Z(NET_628),.Q3Z(m1_ram_control[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_T16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_82),.B0I1(m1_m1_dataout_int[0]),.B0I2(tcdm_result_p2[0]),.B0I3(NET_83),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[6]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T0I0(NET_82),.T0I1(m1_m1_dataout_int[0]),.T0I2(tcdm_result_p2[0]),.T0I3(NET_83),.TB0S(NET_84),.C0Z(NET_80),.Q0Z(tcdm_result_p2[6]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B1I0(tcdm_result_p2[7]),.B1I1(m1_m1_dataout_int[7]),.B1I2(NET_83),.B1I3(NET_82),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T1I0(NET_83),.T1I1(NET_82),.T1I2(tcdm_result_p2[7]),.T1I3(m1_m1_dataout_int[7]),.TB1S(NET_462),.C1Z(NET_460),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_T16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_82),.B2I1(m1_m1_dataout_int[6]),.B2I2(NET_83),.B2I3(tcdm_result_p2[6]),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[0]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T2I0(NET_82),.T2I1(m1_m1_dataout_int[6]),.T2I2(NET_83),.T2I3(tcdm_result_p2[6]),.TB2S(NET_628),.C2Z(NET_626),.Q2Z(tcdm_result_p2[0]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_T16_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[7]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_20_padClk),.QRT(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF),.QST(GND),.T3I0(NET_86),.T3I1(m1_m1_dataout_int[17]),.T3I2(m0_m1_dataout_int[17]),.T3I3(NET_83),.TB3S(GND),.C3Z(NET_335),.Q3Z(tcdm_result_p2[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_T17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m1_m1_dataout_int[12]),.B0I1(NET_83_CAND2_BRSTL_20_tpGCLKBUF),.B0I2(NET_82),.B0I3(tcdm_result_p2[12]),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[14]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.T0I0(m1_m1_dataout_int[12]),.T0I1(NET_83_CAND2_BRSTL_20_tpGCLKBUF),.T0I2(NET_82),.T0I3(tcdm_result_p2[12]),.TB0S(NET_216),.C0Z(NET_214),.Q0Z(tcdm_result_p2[14]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[15]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_T17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[12]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p2[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_U12_0 (.tFragBitInfo(16'b0100110001001100),.bFragBitInfo(16'b0000000001001100),.B0I0(m0_m1_dataout_int[8]),.B0I1(NET_739),.B0I2(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.B0I3(tcdm_result_p1[8]),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[13]),.Q0EN(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T0I0(m0_m1_dataout_int[8]),.T0I1(NET_739),.T0I2(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.T0I3(tcdm_result_p1[8]),.TB0S(NET_50),.C0Z(NET_740),.Q0Z(tcdm_result_p1[13]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[11]),.Q2EN(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p1[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U12_3 (.tFragBitInfo(16'b0100110001001100),.bFragBitInfo(16'b0001001100000000),.B3I0(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.B3I1(tcdm_result_p1[13]),.B3I2(m0_m1_dataout_int[13]),.B3I3(NET_735),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[8]),.Q3EN(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(m0_m1_dataout_int[13]),.T3I1(NET_735),.T3I2(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.T3I3(tcdm_result_p1[13]),.TB3S(NET_50),.C3Z(NET_736),.Q3Z(tcdm_result_p1[8]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_U13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_35),.B0I1(NET_34),.B0I2(tcdm_rdata_p1_int[11]),.B0I3(tcdm_rdata_p3_int[11]),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[9]),.Q0EN(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B0Z(NET_199),.Q0Z(tcdm_result_p1[9]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U13_1 (.tFragBitInfo(16'b0101111100000000),.bFragBitInfo(16'b0000000001001100),.B1I0(m0_m1_dataout_int[10]),.B1I1(NET_731),.B1I2(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.B1I3(tcdm_result_p1[10]),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T1I0(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.T1I1(tcdm_result_p1[10]),.T1I2(m0_m1_dataout_int[10]),.T1I3(NET_731),.TB1S(NET_50),.C1Z(NET_732),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_U13_2 (.tFragBitInfo(16'b0101111100000000),.bFragBitInfo(16'b0001001100000000),.B2I0(m0_m1_dataout_int[9]),.B2I1(tcdm_result_p1[9]),.B2I2(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.B2I3(NET_729),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[10]),.Q2EN(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T2I0(m0_m1_dataout_int[9]),.T2I1(tcdm_result_p1[9]),.T2I2(NET_52_CAND2_TRSBL_21_tpGCLKBUF),.T2I3(NET_729),.TB2S(NET_50),.C2Z(NET_730),.Q2Z(tcdm_result_p1[10]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_U13_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(NET_35),.T3I1(NET_34),.T3I2(tcdm_rdata_p1_int[9]),.T3I3(tcdm_rdata_p3_int[9]),.TB3S(GND),.C3Z(NET_158),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_U14_0 (.tFragBitInfo(16'b0111111101111111),.bFragBitInfo(16'b0000111101111111),.B0I0(NET_49_CAND4_TRSBL_21_tpGCLKBUF),.B0I1(tcdm_result_p3[11]),.B0I2(NET_7_CAND3_TRSBL_21_tpGCLKBUF),.B0I3(tcdm_result_p2[11]),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T0I0(NET_49_CAND4_TRSBL_21_tpGCLKBUF),.T0I1(tcdm_result_p3[11]),.T0I2(NET_7_CAND3_TRSBL_21_tpGCLKBUF),.T0I3(tcdm_result_p2[11]),.TB0S(NET_14),.C0Z(NET_733),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U14_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[11]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p3_int[10]),.T1I1(NET_35),.T1I2(tcdm_rdata_p1_int[10]),.T1I3(NET_34),.C1Z(NET_180),.Q1Z(tcdm_result_p3[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_U14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(tcdm_rdata_p1_int[8]),.B2I1(NET_35),.B2I2(tcdm_rdata_p3_int[8]),.B2I3(NET_34),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[9]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B2Z(NET_279),.Q2Z(tcdm_result_p3[9]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U14_3 (.tFragBitInfo(16'b0101111111111111),.bFragBitInfo(16'b0101010101111111),.B3I0(NET_7_CAND3_TRSBL_21_tpGCLKBUF),.B3I1(NET_49_CAND4_TRSBL_21_tpGCLKBUF),.B3I2(tcdm_result_p3[9]),.B3I3(tcdm_result_p2[9]),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[11]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p3[9]),.T3I1(tcdm_result_p2[9]),.T3I2(NET_7_CAND3_TRSBL_21_tpGCLKBUF),.T3I3(NET_49_CAND4_TRSBL_21_tpGCLKBUF),.TB3S(NET_14),.C3Z(NET_729),.Q3Z(tcdm_result_p2[11]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_U15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[8]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p3[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U15_1 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0000011111111111),.B1I0(tcdm_result_p3[10]),.B1I1(NET_49_CAND4_TRSBL_21_tpGCLKBUF),.B1I2(tcdm_result_p2[10]),.B1I3(NET_7_CAND3_TRSBL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p2[10]),.T1I1(NET_7_CAND3_TRSBL_21_tpGCLKBUF),.T1I2(tcdm_result_p3[10]),.T1I3(NET_49_CAND4_TRSBL_21_tpGCLKBUF),.TB1S(NET_14),.C1Z(NET_731),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_U15_2 (.tFragBitInfo(16'b0111011111111111),.bFragBitInfo(16'b0011011100111111),.B2I0(tcdm_result_p3[8]),.B2I1(NET_7_CAND3_TRSBL_21_tpGCLKBUF),.B2I2(tcdm_result_p2[8]),.B2I3(NET_49_CAND4_TRSBL_21_tpGCLKBUF),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[8]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p3[8]),.T2I1(NET_7_CAND3_TRSBL_21_tpGCLKBUF),.T2I2(tcdm_result_p2[8]),.T2I3(NET_49_CAND4_TRSBL_21_tpGCLKBUF),.TB2S(NET_14),.C2Z(NET_739),.Q2Z(tcdm_result_p2[8]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_U15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[10]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p3[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_U16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[9]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p2[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U16_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[2]),.T3I1(NET_65),.T3I2(GND),.T3I3(GND),.TB3S(GND),.C3Z(NET_145),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_U17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[10]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p2[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V12_0 (.tFragBitInfo(16'b0101000011110000),.bFragBitInfo(16'b0001000000110000),.B0I0(NET_52_CAND2_TRSBL_22_tpGCLKBUF),.B0I1(tcdm_result_p1[3]),.B0I2(NET_760),.B0I3(m0_m1_dataout_int[3]),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[1]),.Q0EN(tcdm_valid_p1_int_CAND5_TRSBL_22_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T0I0(NET_52_CAND2_TRSBL_22_tpGCLKBUF),.T0I1(tcdm_result_p1[3]),.T0I2(NET_760),.T0I3(m0_m1_dataout_int[3]),.TB0S(NET_50),.C0Z(NET_761),.Q0Z(tcdm_result_p1[1]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_V12_1 (.tFragBitInfo(16'b0000110011001100),.bFragBitInfo(16'b0000011100000000),.B1I0(m0_m1_dataout_int[1]),.B1I1(NET_52_CAND2_TRSBL_22_tpGCLKBUF),.B1I2(tcdm_result_p1[1]),.B1I3(NET_727),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p1[1]),.T1I1(NET_727),.T1I2(m0_m1_dataout_int[1]),.T1I3(NET_52_CAND2_TRSBL_22_tpGCLKBUF),.TB1S(NET_50),.C1Z(NET_728),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_V12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[3]),.Q2EN(tcdm_valid_p1_int_CAND5_TRSBL_22_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p1[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V13_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p1_int[3]),.T0I1(NET_35),.T0I2(NET_34),.T0I3(tcdm_rdata_p3_int[3]),.TB0S(GND),.C0Z(NET_692),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_V13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V13_2 (.tFragBitInfo(16'b0111011111111111),.bFragBitInfo(16'b0101011101011111),.B2I0(NET_7_CAND3_TRSBL_22_tpGCLKBUF),.B2I1(NET_49_CAND4_TRSBL_22_tpGCLKBUF),.B2I2(tcdm_result_p2[3]),.B2I3(tcdm_result_p3[3]),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[4]),.Q2EN(tcdm_valid_p1_int_CAND5_TRSBL_22_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T2I0(NET_7_CAND3_TRSBL_22_tpGCLKBUF),.T2I1(NET_49_CAND4_TRSBL_22_tpGCLKBUF),.T2I2(tcdm_result_p2[3]),.T2I3(tcdm_result_p3[3]),.TB2S(NET_14),.C2Z(NET_760),.Q2Z(tcdm_result_p1[4]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_V13_3 (.tFragBitInfo(16'b0000110011001100),.bFragBitInfo(16'b0000011100000000),.B3I0(m0_m1_dataout_int[4]),.B3I1(NET_52_CAND2_TRSBL_22_tpGCLKBUF),.B3I2(tcdm_result_p1[4]),.B3I3(NET_758),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[3]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p1[4]),.T3I1(NET_758),.T3I2(m0_m1_dataout_int[4]),.T3I3(NET_52_CAND2_TRSBL_22_tpGCLKBUF),.TB3S(NET_50),.C3Z(NET_759),.Q3Z(tcdm_result_p3[3]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_V14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_34),.B0I1(NET_35),.B0I2(tcdm_rdata_p1_int[13]),.B0I3(tcdm_rdata_p3_int[13]),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[4]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B0Z(NET_239),.Q0Z(tcdm_result_p3[4]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V14_1 (.tFragBitInfo(16'b0111011111111111),.bFragBitInfo(16'b0011011101110111),.B1I0(tcdm_result_p2[4]),.B1I1(NET_7_CAND3_TRSBL_22_tpGCLKBUF),.B1I2(tcdm_result_p3[4]),.B1I3(NET_49_CAND4_TRSBL_22_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p3[4]),.T1I1(NET_49_CAND4_TRSBL_22_tpGCLKBUF),.T1I2(tcdm_result_p2[4]),.T1I3(NET_7_CAND3_TRSBL_22_tpGCLKBUF),.TB1S(NET_14),.C1Z(NET_758),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_V14_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_34),.B2I1(NET_35),.B2I2(tcdm_rdata_p1_int[1]),.B2I3(tcdm_rdata_p3_int[1]),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T2I0(NET_34),.T2I1(NET_35),.T2I2(tcdm_rdata_p1_int[4]),.T2I3(tcdm_rdata_p3_int[4]),.TB2S(GND),.B2Z(NET_24),.C2Z(NET_673),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_V14_3 (.tFragBitInfo(16'b0111111101111111),.bFragBitInfo(16'b0001111100111111),.B3I0(tcdm_result_p3[1]),.B3I1(tcdm_result_p2[1]),.B3I2(NET_7_CAND3_TRSBL_22_tpGCLKBUF),.B3I3(NET_49_CAND4_TRSBL_22_tpGCLKBUF),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[1]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T3I0(NET_7_CAND3_TRSBL_22_tpGCLKBUF),.T3I1(NET_49_CAND4_TRSBL_22_tpGCLKBUF),.T3I2(tcdm_result_p3[1]),.T3I3(tcdm_result_p2[1]),.TB3S(NET_14),.C3Z(NET_727),.Q3Z(tcdm_result_p3[1]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_V15_0 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0011011101110111),.B0I0(tcdm_result_p2[13]),.B0I1(NET_7_CAND3_TRSBL_22_tpGCLKBUF),.B0I2(NET_49_CAND4_TRSBL_22_tpGCLKBUF),.B0I3(tcdm_result_p3[13]),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p2[13]),.T0I1(NET_7_CAND3_TRSBL_22_tpGCLKBUF),.T0I2(NET_49_CAND4_TRSBL_22_tpGCLKBUF),.T0I3(tcdm_result_p3[13]),.TB0S(NET_14),.C0Z(NET_735),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_V15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[13]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p3[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[4]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p2[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[3]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND1_BRSTL_22_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[1]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND1_BRSTL_22_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND1_BRSTL_22_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[13]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND1_BRSTL_22_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p2[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V18_2 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'b0000000000000000),.T2I0(lint_ADDR_int[4]),.T2I1(lint_ADDR_int[5]),.T2I2(lint_ADDR_int[3]),.T2I3(lint_ADDR_int[6]),.TB2S(GND),.C2Z(NET_7),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_V18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_W3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(NET_762),.Q2EN(nx25587z1),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_we_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_W30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND1_BRSBL_23_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND1_BRSBL_23_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(NET_762),.Q2EN(nx30664z1),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND1_BRSBL_23_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_we_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND1_BRSBL_23_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx25587z1),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[11]),.Q1EN(nx25587z1),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_waddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[11]),.Q2EN(nx18281z1),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_raddr_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx25587z1),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx30664z1),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND1_BRSBL_24_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[11]),.Q1EN(nx53672z1),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND1_BRSBL_24_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_raddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND1_BRSBL_24_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[11]),.Q3EN(nx30664z1),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND1_BRSBL_24_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_waddr_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx30664z1),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND1_BRSBL_24_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND1_BRSBL_24_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND1_BRSBL_24_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx30664z1),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND1_BRSBL_24_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[29]),.Q0EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[29]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[23]),.Q2EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[21]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[20]),.Q2EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[20]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y19_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_65),.T2I1(GND),.T2I2(GND),.T2I3(NET_134),.TB2S(GND),.C2Z(NET_133),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_Y19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[20]),.Q2EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[20]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[19]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[6]),.Q2EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_waddr_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_wdata_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_wdata_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wdata_dup_0[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z17_2 (.tFragBitInfo(16'b0000000000000100),.bFragBitInfo(16'b0000010000000000),.B2I0(GND),.B2I1(NET_65),.B2I2(GND),.B2I3(lint_ADDR_int[3]),.T2I0(lint_ADDR_int[2]),.T2I1(NET_65),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(NET_645),.C2Z(NET_135),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_Z17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_wdata_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_wdata_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[3]),.Q1EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_waddr_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_wdata_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[9]),.Q3EN(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_waddr_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[0]),.Q0EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_waddr_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[9]),.Q1EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_waddr_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[5]),.Q2EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_waddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_waddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[7]),.Q0EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_waddr_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[4]),.Q1EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_waddr_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[2]),.Q2EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_waddr_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[1]),.Q3EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_waddr_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[3]),.Q1EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_waddr_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[8]),.Q2EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_waddr_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdata_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(lint_ADDR_int[3]),.B0I1(GND),.B0I2(GND),.B0I3(lint_ADDR_int[2]),.B0Z(NET_138),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[6]),.Q2EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_waddr_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_wdata_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[5]),.Q0EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_waddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[10]),.Q1EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_waddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[2]),.Q2EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_waddr_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[4]),.Q3EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_waddr_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[7]),.Q0EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_waddr_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[0]),.Q1EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_waddr_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[8]),.Q2EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_waddr_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[1]),.Q3EN(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_waddr_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[4]),.Q0EN(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_raddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[10]),.Q1EN(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_raddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[6]),.Q2EN(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_raddr_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[5]),.Q3EN(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_raddr_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[8]),.Q1EN(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_raddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[3]),.Q2EN(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_raddr_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB8_1 (.tFragBitInfo(16'b1111000011110000),.bFragBitInfo(16'b1110101010101010),.B1I0(tcdm_gnt_p0_int),.B1I1(NET_65),.B1I2(NET_131),.B1I3(NET_138),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.T1I0(NET_131),.T1I1(NET_138),.T1I2(tcdm_gnt_p0_int),.T1I3(NET_65),.TB1S(NET_132),.C1Z(nx11313z3),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_AB8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_172),.B2I1(NET_138),.B2I2(NET_132),.B2I3(NET_65),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.T2I0(NET_172),.T2I1(NET_138),.T2I2(NET_132),.T2I3(NET_65),.TB2S(lint_ADDR_int[7]),.C2Z(nx41193z1),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_AB8_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx11313z3),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.T3I0(NET_132),.T3I1(NET_138),.T3I2(NET_65),.T3I3(NET_131),.TB3S(GND),.Q3Z(tcdm_req_p0_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB9_1 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[2]),.T1I1(lint_ADDR_int[3]),.T1I2(GND),.T1I3(NET_65),.C1Z(NET_137),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_AB9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B0I0(lint_ADDR_int[2]),.B0I1(lint_ADDR_int[3]),.B0I2(GND),.B0I3(lint_ADDR_int[7]),.B0Z(NET_386),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB11_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_65),.T1I1(NET_386),.T1I2(NET_172),.T1I3(NET_132),.TB1S(GND),.C1Z(nx36058z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_AB11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB11_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int[5]),.T3I1(lint_ADDR_int[4]),.T3I2(GND),.T3I3(GND),.C3Z(NET_172),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_AB17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND1_BRSTR_28_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB17_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx11311z2),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND1_BRSTR_28_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[3]),.T1I1(NET_135),.T1I2(NET_131),.T1I3(NET_132),.TB1S(GND),.Q1Z(tcdm_req_p2_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AB17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1111111110000000),.B2I0(NET_131),.B2I1(NET_132),.B2I2(NET_136),.B2I3(tcdm_gnt_p2_int),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND1_BRSTR_28_tpGCLKBUF),.QST(GND),.B2Z(nx11311z2),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB17_3 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND1_BRSTR_28_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[3]),.T3I1(GND),.T3I2(lint_ADDR_int[2]),.T3I3(NET_65),.C3Z(NET_136),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_AB18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB18_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int[7]),.T3I1(lint_ADDR_int[4]),.T3I2(lint_ADDR_int[5]),.T3I3(GND),.C3Z(NET_131),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_AB19_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.T0I0(NET_134),.T0I1(RESET_int[0]),.T0I2(NET_172),.T0I3(NET_65),.TB0S(GND),.C0Z(NET_666),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_AB19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB19_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000001000000000),.B2I0(lint_ADDR_int[3]),.B2I1(lint_ADDR_int[2]),.B2I2(GND),.B2I3(lint_ADDR_int[7]),.T2I0(NET_132),.T2I1(NET_272),.T2I2(NET_172),.T2I3(NET_65),.TB2S(GND),.B2Z(NET_272),.C2Z(nx30923z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_AB19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_65),.B0I1(NET_134),.B0I2(NET_132),.B0I3(NET_172),.T0I0(NET_65),.T0I1(NET_134),.T0I2(NET_132),.T0I3(NET_172),.TB0S(lint_ADDR_int[7]),.C0Z(nx25788z1),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_AB20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[6]),.Q0EN(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_raddr_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[4]),.Q1EN(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_raddr_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[5]),.Q2EN(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_raddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[10]),.Q1EN(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_raddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[3]),.Q2EN(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_raddr_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[8]),.Q3EN(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_raddr_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[0]),.Q0EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q0Z(m0_oper1_raddr_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[1]),.Q1EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper1_raddr_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[9]),.Q2EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_raddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[2]),.Q2EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_raddr_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[7]),.Q3EN(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_raddr_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx41193z1_CAND3_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[21]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1110101010101010),.B0I0(tcdm_gnt_p1_int),.B0I1(NET_132),.B0I2(NET_137),.B0I3(NET_131),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B0Z(nx11312z2),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC9_3 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx11312z2),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_132),.T3I2(NET_137),.T3I3(NET_131),.TB3S(GND),.Q3Z(tcdm_req_p1_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AC10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[8]),.Q1EN(nx52746z1_CAND3_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx36058z1_CAND2_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx52746z1_CAND3_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p1_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[8]),.Q1EN(nx36058z1_CAND2_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx36058z1_CAND2_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[21]),.Q1EN(nx36058z1_CAND2_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC14_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_145),.T1I1(NET_147),.T1I2(RESET_int[0]),.T1I3(NET_146),.TB1S(GND),.C1Z(nx16907z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_AC14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC14_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_145),.T3I1(NET_147),.T3I2(NET_146),.T3I3(GND),.TB3S(GND),.C3Z(nx52746z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_AC20_0 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000010000000),.B0I0(NET_147),.B0I1(NET_666),.B0I2(NET_132),.B0I3(GND),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.T0I0(NET_147),.T0I1(NET_133),.T0I2(NET_132),.T0I3(GND),.TB0S(GND),.B0Z(nx65467z1),.C0Z(nx2520z1),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AC20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC20_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx11310z2),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.T2I0(NET_131),.T2I1(NET_133),.T2I2(NET_132),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_req_p3_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AC20_3 (.tFragBitInfo(16'b1111111110000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[21]),.Q3EN(nx30923z1_CAND4_BRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF),.QST(GND),.T3I0(NET_131),.T3I1(NET_133),.T3I2(NET_132),.T3I3(tcdm_gnt_p3_int),.C3Z(nx11310z2),.Q3Z(tcdm_wdata_p2_dup_0[21]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_AC26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx25788z1_CAND3_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[2]),.Q1EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_raddr_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[7]),.Q0EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q0Z(m1_oper1_raddr_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[1]),.Q1EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q1Z(m1_oper1_raddr_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[0]),.Q2EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_raddr_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[9]),.Q3EN(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper1_raddr_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx47611z1_CAND4_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p0_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx47611z1_CAND4_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p0_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[20]),.Q3EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_30_padClk),.QRT(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_BE_int[3]),.Q0EN(nx16907z1),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_be_p1_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_BE_int[0]),.Q1EN(nx16907z1),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_be_p1_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_BE_int[0]),.Q2EN(nx25326z1),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_be_p0_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_BE_int[3]),.Q3EN(nx25326z1),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_be_p0_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx52746z1_CAND3_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p1_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_BE_int[2]),.Q0EN(nx25326z1),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_be_p0_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_BE_int[2]),.Q2EN(nx16907z1),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_be_p1_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(GND),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx52746z1_CAND3_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_30_padClk),.QRT(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD14_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_147),.T1I1(NET_173),.T1I2(GND),.T1I3(NET_68),.C1Z(nx47611z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_AD14_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_147),.T2I1(NET_173),.T2I2(RESET_int[0]),.T2I3(NET_68),.TB2S(GND),.C2Z(nx25326z1),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_AD14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD16_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_147),.T1I1(NET_68),.T1I2(GND),.T1I3(NET_645),.C1Z(nx57881z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_AD16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_BE_int[0]),.Q0EN(nx8488z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_be_p2_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_BE_int[2]),.Q1EN(nx8488z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_be_p2_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD17_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_BE_int[3]),.Q3EN(nx8488z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.T3I0(RESET_int[0]),.T3I1(NET_68),.T3I2(NET_645),.T3I3(NET_147),.TB3S(GND),.C3Z(nx8488z1),.Q3Z(tcdm_be_p2_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_AD18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx57881z1_CAND3_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p2_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx57881z1_CAND3_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[9]),.Q1EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx57881z1_CAND3_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[23]),.Q1EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[23]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_BE_int[3]),.Q0EN(nx65467z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_be_p3_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx65467z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_we_p3_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_BE_int[2]),.Q1EN(nx65467z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_be_p3_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_BE_int[1]),.Q2EN(nx65467z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_be_p3_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_BE_int[0]),.Q3EN(nx65467z1),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_be_p3_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx2520z1_CAND2_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p3_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx2520z1_CAND2_BRSTR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_30_padClk),.QRT(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx2520z1_CAND2_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p3_dup_0[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AD27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AD27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AD27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[30]),.Q2EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[30]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AD27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_30_padClk),.QRT(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p0_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p0_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p0_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p0_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[18]),.Q2EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[18]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_31_padClk),.QRT(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_BE_int[1]),.Q0EN(nx25326z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_be_p0_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx16907z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_we_p1_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_BE_int[1]),.Q2EN(nx16907z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_be_p1_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx25326z1),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_we_p0_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p1_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p1_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[17]),.Q0EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[17]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p1_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p1_dup_0[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_31_padClk),.QRT(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(GND),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(GND),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx8488z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_we_p2_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_BE_int[1]),.Q3EN(nx8488z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_be_p2_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p2_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p2_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p2_dup_0[13]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p2_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[18]),.Q2EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[18]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p2_dup_0[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx2520z1_CAND2_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p3_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx2520z1_CAND2_BRSTR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_31_padClk),.QRT(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[13]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p3_dup_0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p3_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p3_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[14]),.Q3EN(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p3_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AE27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[25]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AE27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p3_dup_0[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AE27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AE27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[24]),.Q3EN(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_31_padClk),.QRT(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p0_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p0_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[17]),.Q0EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p0_dup_0[17]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p0_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p0_dup_0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[26]),.Q1EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p0_dup_0[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p0_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_32_padClk),.QRT(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p0_dup_0[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p1_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p1_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p1_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p1_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p1_dup_0[12]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[9]),.Q1EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p1_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p1_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p1_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p1_dup_0[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p1_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p1_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p1_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx57881z1),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p2_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx57881z1),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_32_padClk),.QRT(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p2_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p2_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p2_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p2_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p2_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p2_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p2_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p2_dup_0[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p2_dup_0[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p2_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p2_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p2_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p3_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_addr_p3_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p3_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx25788z1),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_32_padClk),.QRT(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p3_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx2520z1_CAND2_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p3_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p3_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx2520z1_CAND2_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p3_dup_0[19]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx2520z1_CAND2_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AF27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[28]),.Q0EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_wdata_p3_dup_0[28]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AF27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_wdata_p3_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AF27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_wdata_p3_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AF27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_32_padClk),.QRT(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_wdata_p3_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	CLOCK QL_INST_IO_CLK0 (.CEN(VCC),.IP(CLK[0]),.IC(CLK_int[0]),.OP());

	CLOCK QL_INST_IO_CLK1 (.CEN(VCC),.IP(CLK[1]),.IC(CLK_int[1]),.OP());

	CLOCK QL_INST_IO_CLK2 (.CEN(VCC),.IP(CLK[2]),.IC(CLK_int[2]),.OP());

	CLOCK QL_INST_IO_CLK3 (.CEN(VCC),.IP(CLK[3]),.IC(CLK_int[3]),.OP());

	CLOCK QL_INST_IO_CLK4 (.CEN(VCC),.IP(CLK[4]),.IC(CLK_int[4]),.OP());

	CLOCK QL_INST_IO_CLK5 (.CEN(VCC),.IP(CLK[5]),.IC(CLK_int[5]),.OP());

	GMUX QL_INST_GMUX_0 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[0]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_0__GMUX_0_padClk));

	GMUX QL_INST_GMUX_1 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[1]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_1__GMUX_1_padClk));

	GMUX QL_INST_GMUX_2 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[2]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_2__GMUX_2_padClk));

	GMUX QL_INST_GMUX_3 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[3]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_3__GMUX_3_padClk));

	GMUX QL_INST_GMUX_4 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[4]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_4__GMUX_4_padClk));

	GMUX QL_INST_GMUX_5 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[5]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_5__GMUX_5_padClk));

	QPMUX QL_INST_QMUX_TL0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_TL0_padClk));

	QPMUX QL_INST_QMUX_TL1 (.GMUXIN(CLK_int_1__GMUX_1_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_1__QMUX_TL1_padClk));

	QPMUX QL_INST_QMUX_TL2 (.GMUXIN(CLK_int_2__GMUX_2_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_2__QMUX_TL2_padClk));

	QMUX QL_INST_QMUX_TL3 (.GMUXIN(GND),.IS(VCC),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_TL3_tpGCLKBUF));

	QMUX QL_INST_QMUX_TL4 (.GMUXIN(CLK_int_4__GMUX_4_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_4__QMUX_TL4_padClk));

	QMUX QL_INST_QMUX_TL5 (.GMUXIN(CLK_int_5__GMUX_5_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_5__QMUX_TL5_padClk));

	QPMUX QL_INST_QMUX_TR0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_TR0_padClk));

	QPMUX QL_INST_QMUX_TR1 (.GMUXIN(GND),.IS0(VCC),.IS1(VCC),.QCLKIN(GND),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_TR1_tpGCLKBUF));

	QMUX QL_INST_QMUX_BL0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_BL0_padClk));

	QMUX QL_INST_QMUX_BL1 (.GMUXIN(GND),.IS(VCC),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_BL1_tpGCLKBUF));

	QMUX QL_INST_QMUX_BL2 (.GMUXIN(GND),.IS(VCC),.QHSCK(nx9707z1),.IZ(nx9707z1_QMUX_BL2_tpGCLKBUF));

	QPMUX QL_INST_QMUX_BL3 (.GMUXIN(CLK_int_3__GMUX_3_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_3__QMUX_BL3_padClk));

	QMUX QL_INST_QMUX_BR0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_BR0_padClk));

	QMUX QL_INST_QMUX_BR1 (.GMUXIN(GND),.IS(VCC),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_BR1_tpGCLKBUF));

	QMUX QL_INST_QMUX_BR2 (.GMUXIN(GND),.IS(VCC),.QHSCK(nx2520z1),.IZ(nx2520z1_QMUX_BR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSTL0_padClk));

	SQEMUX QL_INST_SQMUX_TLSTL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx44608z1),.IZ(nx44608z1_SQMUX_TLSTL1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx34006z2),.IZ(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTL3 (.QMUXIN(not_RESET_0_QMUX_TL3_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TLSTL3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTL4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx39840z1),.IZ(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTL5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx34850z1),.IZ(nx34850z1_SQMUX_TLSTL5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSTR0_padClk));

	SQEMUX QL_INST_SQMUX_TLSTR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_46),.IZ(NET_46_SQMUX_TLSTR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx15998z1),.IZ(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTR3 (.QMUXIN(not_RESET_0_QMUX_TL3_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TLSTR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTR4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(lint_ADDR_int[13]),.IZ(lint_ADDR_int_13__SQMUX_TLSTR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTR5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(lint_ADDR_int[14]),.IZ(lint_ADDR_int_14__SQMUX_TLSTR5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSBL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSBL0_padClk));

	SQEMUX QL_INST_SQMUX_TLSBL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_1__QMUX_TL1_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_1__SQMUX_TLSBL1_padClk));

	SQEMUX QL_INST_SQMUX_TLSBL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_2__QMUX_TL2_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_2__SQMUX_TLSBL2_padClk));

	SQMUX QL_INST_SQMUX_TLSBL3 (.QMUXIN(not_RESET_0_QMUX_TL3_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TLSBL3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBL4 (.QMUXIN(CLK_int_4__QMUX_TL4_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_4__SQMUX_TLSBL4_padClk));

	SQMUX QL_INST_SQMUX_TLSBL5 (.QMUXIN(CLK_int_5__QMUX_TL5_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_5__SQMUX_TLSBL5_padClk));

	SQEMUX QL_INST_SQMUX_TLSBR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSBR0_padClk));

	SQEMUX QL_INST_SQMUX_TLSBR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(tcdm_valid_p0_int),.IZ(tcdm_valid_p0_int_SQMUX_TLSBR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSBR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx49808z64),.IZ(nx49808z64_SQMUX_TLSBR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBR3 (.QMUXIN(not_RESET_0_QMUX_TL3_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TLSBR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBR4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_124),.IZ(NET_124_SQMUX_TLSBR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBR5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_15),.IZ(NET_15_SQMUX_TLSBR5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSTL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSTL0_padClk));

	SQEMUX QL_INST_SQMUX_TRSTL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSTL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx32231z1),.IZ(nx32231z1_SQMUX_TRSTL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSTR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSTR0_padClk));

	SQEMUX QL_INST_SQMUX_TRSTR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSTR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx25587z1),.IZ(nx25587z1_SQMUX_TRSTR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTR3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx41193z1),.IZ(nx41193z1_SQMUX_TRSTR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTR4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx47611z1),.IZ(nx47611z1_SQMUX_TRSTR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTR5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx18281z1),.IZ(nx18281z1_SQMUX_TRSTR5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSBL0_padClk));

	SQEMUX QL_INST_SQMUX_TRSBL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_52),.IZ(NET_52_SQMUX_TRSBL2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBL3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_7),.IZ(NET_7_SQMUX_TRSBL3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBL4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_49),.IZ(NET_49_SQMUX_TRSBL4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBL5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(tcdm_valid_p1_int),.IZ(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSBR0_padClk));

	SQEMUX QL_INST_SQMUX_TRSBR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx36058z1),.IZ(nx36058z1_SQMUX_TRSBR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBR3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx52746z1),.IZ(nx52746z1_SQMUX_TRSBR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTL0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSTL0_padClk));

	SQMUX QL_INST_SQMUX_BLSTL1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTL2 (.QMUXIN(nx9707z1_QMUX_BL2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTL3 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_3__QMUX_BL3_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_3__SQMUX_BLSTL3_padClk));

	SQEMUX QL_INST_SQMUX_BLSTL4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx4939z1),.IZ(nx4939z1_SQMUX_BLSTL4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTL5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_29),.IZ(NET_29_SQMUX_BLSTL5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTR0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSTR0_padClk));

	SQMUX QL_INST_SQMUX_BLSTR1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTR2 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx19726z1),.IZ(nx19726z1_SQMUX_BLSTR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_17),.IZ(NET_17_SQMUX_BLSTR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_28),.IZ(NET_28_SQMUX_BLSTR4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTR5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_18),.IZ(NET_18_SQMUX_BLSTR5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBL0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSBL0_padClk));

	SQMUX QL_INST_SQMUX_BLSBL1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBL2 (.QMUXIN(nx9707z1_QMUX_BL2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBL3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx60831z1),.IZ(nx60831z1_SQMUX_BLSBL3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBL4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx22245z1),.IZ(nx22245z1_SQMUX_BLSBL4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBR0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSBR0_padClk));

	SQMUX QL_INST_SQMUX_BLSBR1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBR2 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx33579z1),.IZ(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_43),.IZ(NET_43_SQMUX_BLSBR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_44),.IZ(NET_44_SQMUX_BLSBR4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBR5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_32),.IZ(NET_32_SQMUX_BLSBR5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTL0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSTL0_padClk));

	SQMUX QL_INST_SQMUX_BRSTL1 (.QMUXIN(not_RESET_0_QMUX_BR1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTL2 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_83),.IZ(NET_83_SQMUX_BRSTL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTL3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_125),.IZ(NET_125_SQMUX_BRSTL3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTL4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_110),.IZ(NET_110_SQMUX_BRSTL4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTR0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSTR0_padClk));

	SQMUX QL_INST_SQMUX_BRSTR1 (.QMUXIN(not_RESET_0_QMUX_BR1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTR2 (.QMUXIN(nx2520z1_QMUX_BR2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(nx2520z1_SQMUX_BRSTR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx57881z1),.IZ(nx57881z1_SQMUX_BRSTR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx30923z1),.IZ(nx30923z1_SQMUX_BRSTR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSBL0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSBL0_padClk));

	SQMUX QL_INST_SQMUX_BRSBL1 (.QMUXIN(not_RESET_0_QMUX_BR1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSBL1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSBL2 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx14650z1),.IZ(nx14650z1_SQMUX_BRSBL2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSBR0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSBR0_padClk));

	SQMUX QL_INST_SQMUX_BRSBR1 (.QMUXIN(not_RESET_0_QMUX_BR1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSBR2 (.QMUXIN(nx2520z1_QMUX_BR2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(nx2520z1_SQMUX_BRSBR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx25788z1),.IZ(nx25788z1_SQMUX_BRSBR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx53672z1),.IZ(nx53672z1_SQMUX_BRSBR4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBR5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx30664z1),.IZ(nx30664z1_SQMUX_BRSBR5_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSTL_1 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_1_padClk));

	CAND QL_INST_CAND0_TLSTL_2 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_2_padClk));

	CAND QL_INST_CAND0_TLSTL_3 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_3_padClk));

	CAND QL_INST_CAND0_TLSTL_4 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_4_padClk));

	CAND QL_INST_CAND0_TLSTL_5 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_5_padClk));

	CAND QL_INST_CAND0_TLSTL_6 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_6_padClk));

	CAND QL_INST_CAND0_TLSTL_7 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_7_padClk));

	CAND QL_INST_CAND0_TLSTL_8 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_8_padClk));

	CAND QL_INST_CAND1_TLSTL_1 (.CLKIN(nx44608z1_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(nx44608z1_CAND1_TLSTL_1_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_2 (.CLKIN(nx44608z1_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(nx44608z1_CAND1_TLSTL_2_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_3 (.CLKIN(nx44608z1_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(nx44608z1_CAND1_TLSTL_3_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_5 (.CLKIN(nx44608z1_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(nx44608z1_CAND1_TLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_4 (.CLKIN(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_5 (.CLKIN(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_6 (.CLKIN(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_7 (.CLKIN(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z2_CAND2_TLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_1 (.CLKIN(not_RESET_0_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_2 (.CLKIN(not_RESET_0_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_3 (.CLKIN(not_RESET_0_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_4 (.CLKIN(not_RESET_0_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_5 (.CLKIN(not_RESET_0_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_6 (.CLKIN(not_RESET_0_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_7 (.CLKIN(not_RESET_0_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_8 (.CLKIN(not_RESET_0_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_3 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_4 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_5 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_6 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_7 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_8 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTL_7 (.CLKIN(nx34850z1_SQMUX_TLSTL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx34850z1_CAND5_TLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTL_8 (.CLKIN(nx34850z1_SQMUX_TLSTL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx34850z1_CAND5_TLSTL_8_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSTR_9 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_9_padClk));

	CAND QL_INST_CAND0_TLSTR_12 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_12_padClk));

	CAND QL_INST_CAND0_TLSTR_13 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_13_padClk));

	CAND QL_INST_CAND0_TLSTR_14 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_14_padClk));

	CAND QL_INST_CAND0_TLSTR_15 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_15_padClk));

	CAND QL_INST_CAND0_TLSTR_16 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_16_padClk));

	CAND QL_INST_CAND1_TLSTR_11 (.CLKIN(NET_46_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(NET_46_CAND1_TLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_12 (.CLKIN(NET_46_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(NET_46_CAND1_TLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_13 (.CLKIN(NET_46_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(NET_46_CAND1_TLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_14 (.CLKIN(NET_46_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(NET_46_CAND1_TLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_15 (.CLKIN(NET_46_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(NET_46_CAND1_TLSTR_15_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_16 (.CLKIN(NET_46_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(NET_46_CAND1_TLSTR_16_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_13 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_14 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_15 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_15_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_16 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_9 (.CLKIN(not_RESET_0_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_12 (.CLKIN(not_RESET_0_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_13 (.CLKIN(not_RESET_0_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_14 (.CLKIN(not_RESET_0_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_15 (.CLKIN(not_RESET_0_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_16 (.CLKIN(not_RESET_0_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSTR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_10 (.CLKIN(lint_ADDR_int_13__SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_13__CAND4_TLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_11 (.CLKIN(lint_ADDR_int_13__SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_13__CAND4_TLSTR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_12 (.CLKIN(lint_ADDR_int_13__SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_13__CAND4_TLSTR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_13 (.CLKIN(lint_ADDR_int_13__SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_13__CAND4_TLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_14 (.CLKIN(lint_ADDR_int_13__SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_13__CAND4_TLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_15 (.CLKIN(lint_ADDR_int_13__SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_13__CAND4_TLSTR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTR_10 (.CLKIN(lint_ADDR_int_14__SQMUX_TLSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_14__CAND5_TLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTR_11 (.CLKIN(lint_ADDR_int_14__SQMUX_TLSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_14__CAND5_TLSTR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTR_12 (.CLKIN(lint_ADDR_int_14__SQMUX_TLSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_14__CAND5_TLSTR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTR_13 (.CLKIN(lint_ADDR_int_14__SQMUX_TLSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_14__CAND5_TLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTR_14 (.CLKIN(lint_ADDR_int_14__SQMUX_TLSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_14__CAND5_TLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSBL_1 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_1_padClk));

	CAND QL_INST_CAND0_TLSBL_3 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_3_padClk));

	CAND QL_INST_CAND0_TLSBL_4 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_4_padClk));

	CAND QL_INST_CAND0_TLSBL_5 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_5_padClk));

	CAND QL_INST_CAND0_TLSBL_6 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_6_padClk));

	CAND QL_INST_CAND0_TLSBL_7 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_7_padClk));

	CAND QL_INST_CAND0_TLSBL_8 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_8_padClk));

	CAND QL_INST_CAND1_TLSBL_8 (.CLKIN(CLK_int_1__SQMUX_TLSBL1_padClk),.SEN(VCC),.IZ(CLK_int_1__CAND1_TLSBL_8_padClk));

	CAND QL_INST_CAND2_TLSBL_8 (.CLKIN(CLK_int_2__SQMUX_TLSBL2_padClk),.SEN(VCC),.IZ(CLK_int_2__CAND2_TLSBL_8_padClk));

	CANDEN QL_INST_CAND3_TLSBL_1 (.CLKIN(not_RESET_0_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_3 (.CLKIN(not_RESET_0_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_4 (.CLKIN(not_RESET_0_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_5 (.CLKIN(not_RESET_0_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_6 (.CLKIN(not_RESET_0_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_7 (.CLKIN(not_RESET_0_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_8 (.CLKIN(not_RESET_0_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBL_8 (.CLKIN(CLK_int_4__SQMUX_TLSBL4_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_4__CAND4_TLSBL_8_padClk));

	CANDEN QL_INST_CAND5_TLSBL_7 (.CLKIN(CLK_int_5__SQMUX_TLSBL5_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_5__CAND5_TLSBL_7_padClk));

	CAND QL_INST_CAND0_TLSBR_9 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_9_padClk));

	CAND QL_INST_CAND0_TLSBR_10 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_10_padClk));

	CAND QL_INST_CAND0_TLSBR_11 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_11_padClk));

	CAND QL_INST_CAND0_TLSBR_12 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_12_padClk));

	CAND QL_INST_CAND0_TLSBR_13 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_13_padClk));

	CAND QL_INST_CAND0_TLSBR_14 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_14_padClk));

	CAND QL_INST_CAND0_TLSBR_15 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_15_padClk));

	CAND QL_INST_CAND0_TLSBR_16 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_16_padClk));

	CAND QL_INST_CAND1_TLSBR_12 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND1_TLSBR_12_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_13 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND1_TLSBR_13_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_14 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND1_TLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_15 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND1_TLSBR_15_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_16 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND1_TLSBR_16_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_9 (.CLKIN(nx49808z64_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx49808z64_CAND2_TLSBR_9_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_10 (.CLKIN(nx49808z64_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx49808z64_CAND2_TLSBR_10_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_11 (.CLKIN(nx49808z64_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx49808z64_CAND2_TLSBR_11_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_12 (.CLKIN(nx49808z64_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx49808z64_CAND2_TLSBR_12_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_13 (.CLKIN(nx49808z64_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx49808z64_CAND2_TLSBR_13_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_14 (.CLKIN(nx49808z64_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx49808z64_CAND2_TLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_9 (.CLKIN(not_RESET_0_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_10 (.CLKIN(not_RESET_0_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_11 (.CLKIN(not_RESET_0_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_12 (.CLKIN(not_RESET_0_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_13 (.CLKIN(not_RESET_0_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_14 (.CLKIN(not_RESET_0_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_15 (.CLKIN(not_RESET_0_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_16 (.CLKIN(not_RESET_0_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND3_TLSBR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_12 (.CLKIN(NET_124_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_124_CAND4_TLSBR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_13 (.CLKIN(NET_124_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_124_CAND4_TLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_14 (.CLKIN(NET_124_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_124_CAND4_TLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBR_12 (.CLKIN(NET_15_SQMUX_TLSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_15_CAND5_TLSBR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBR_13 (.CLKIN(NET_15_SQMUX_TLSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_15_CAND5_TLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBR_14 (.CLKIN(NET_15_SQMUX_TLSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_15_CAND5_TLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBR_15 (.CLKIN(NET_15_SQMUX_TLSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_15_CAND5_TLSBR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBR_16 (.CLKIN(NET_15_SQMUX_TLSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_15_CAND5_TLSBR_16_tpGCLKBUF));

	CAND QL_INST_CAND0_TRSTL_17 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_17_padClk));

	CAND QL_INST_CAND0_TRSTL_18 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_18_padClk));

	CAND QL_INST_CAND0_TRSTL_19 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_19_padClk));

	CAND QL_INST_CAND0_TRSTL_23 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_23_padClk));

	CAND QL_INST_CAND0_TRSTL_24 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_24_padClk));

	CAND QL_INST_CAND1_TRSTL_17 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTL_18 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTL_23 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTL_24 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTL_17 (.CLKIN(nx32231z1_SQMUX_TRSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx32231z1_CAND2_TRSTL_17_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTL_18 (.CLKIN(nx32231z1_SQMUX_TRSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx32231z1_CAND2_TRSTL_18_tpGCLKBUF));

	CAND QL_INST_CAND0_TRSTR_25 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_25_padClk));

	CAND QL_INST_CAND0_TRSTR_26 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_26_padClk));

	CAND QL_INST_CAND0_TRSTR_27 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_27_padClk));

	CAND QL_INST_CAND0_TRSTR_28 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_28_padClk));

	CAND QL_INST_CAND0_TRSTR_29 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_29_padClk));

	CAND QL_INST_CAND0_TRSTR_30 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_30_padClk));

	CAND QL_INST_CAND0_TRSTR_31 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_31_padClk));

	CAND QL_INST_CAND0_TRSTR_32 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_32_padClk));

	CAND QL_INST_CAND0_TRSTR_33 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_33_padClk));

	CAND QL_INST_CAND1_TRSTR_25 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_26 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_27 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_28 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_29 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_30 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_30_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_31 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_31_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_32 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_32_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTR_25 (.CLKIN(nx25587z1_SQMUX_TRSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx25587z1_CAND2_TRSTR_25_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTR_26 (.CLKIN(nx25587z1_SQMUX_TRSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx25587z1_CAND2_TRSTR_26_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTR_27 (.CLKIN(nx25587z1_SQMUX_TRSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx25587z1_CAND2_TRSTR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_29 (.CLKIN(nx41193z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z1_CAND3_TRSTR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_30 (.CLKIN(nx41193z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z1_CAND3_TRSTR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_31 (.CLKIN(nx41193z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z1_CAND3_TRSTR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_32 (.CLKIN(nx41193z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z1_CAND3_TRSTR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_30 (.CLKIN(nx47611z1_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx47611z1_CAND4_TRSTR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_31 (.CLKIN(nx47611z1_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx47611z1_CAND4_TRSTR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_32 (.CLKIN(nx47611z1_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx47611z1_CAND4_TRSTR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSTR_28 (.CLKIN(nx18281z1_SQMUX_TRSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx18281z1_CAND5_TRSTR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSTR_29 (.CLKIN(nx18281z1_SQMUX_TRSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx18281z1_CAND5_TRSTR_29_tpGCLKBUF));

	CAND QL_INST_CAND0_TRSBL_17 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_17_padClk));

	CAND QL_INST_CAND0_TRSBL_18 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_18_padClk));

	CAND QL_INST_CAND0_TRSBL_19 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_19_padClk));

	CAND QL_INST_CAND0_TRSBL_20 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_20_padClk));

	CAND QL_INST_CAND0_TRSBL_21 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_21_padClk));

	CAND QL_INST_CAND0_TRSBL_22 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_22_padClk));

	CAND QL_INST_CAND1_TRSBL_17 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_18 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_19 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_20 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_20_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_21 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_22 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBL_18 (.CLKIN(NET_52_SQMUX_TRSBL2_tpGCLKBUF),.SEN(VCC),.IZ(NET_52_CAND2_TRSBL_18_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBL_19 (.CLKIN(NET_52_SQMUX_TRSBL2_tpGCLKBUF),.SEN(VCC),.IZ(NET_52_CAND2_TRSBL_19_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBL_20 (.CLKIN(NET_52_SQMUX_TRSBL2_tpGCLKBUF),.SEN(VCC),.IZ(NET_52_CAND2_TRSBL_20_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBL_21 (.CLKIN(NET_52_SQMUX_TRSBL2_tpGCLKBUF),.SEN(VCC),.IZ(NET_52_CAND2_TRSBL_21_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBL_22 (.CLKIN(NET_52_SQMUX_TRSBL2_tpGCLKBUF),.SEN(VCC),.IZ(NET_52_CAND2_TRSBL_22_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBL_17 (.CLKIN(NET_7_SQMUX_TRSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_7_CAND3_TRSBL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBL_18 (.CLKIN(NET_7_SQMUX_TRSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_7_CAND3_TRSBL_18_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBL_19 (.CLKIN(NET_7_SQMUX_TRSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_7_CAND3_TRSBL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBL_20 (.CLKIN(NET_7_SQMUX_TRSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_7_CAND3_TRSBL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBL_21 (.CLKIN(NET_7_SQMUX_TRSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_7_CAND3_TRSBL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBL_22 (.CLKIN(NET_7_SQMUX_TRSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_7_CAND3_TRSBL_22_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBL_17 (.CLKIN(NET_49_SQMUX_TRSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_49_CAND4_TRSBL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBL_19 (.CLKIN(NET_49_SQMUX_TRSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_49_CAND4_TRSBL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBL_20 (.CLKIN(NET_49_SQMUX_TRSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_49_CAND4_TRSBL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBL_21 (.CLKIN(NET_49_SQMUX_TRSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_49_CAND4_TRSBL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBL_22 (.CLKIN(NET_49_SQMUX_TRSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_49_CAND4_TRSBL_22_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBL_17 (.CLKIN(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p1_int_CAND5_TRSBL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBL_18 (.CLKIN(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p1_int_CAND5_TRSBL_18_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBL_19 (.CLKIN(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p1_int_CAND5_TRSBL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBL_20 (.CLKIN(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p1_int_CAND5_TRSBL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBL_21 (.CLKIN(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p1_int_CAND5_TRSBL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBL_22 (.CLKIN(tcdm_valid_p1_int_SQMUX_TRSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p1_int_CAND5_TRSBL_22_tpGCLKBUF));

	CAND QL_INST_CAND0_TRSBR_29 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_29_padClk));

	CAND QL_INST_CAND0_TRSBR_30 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_30_padClk));

	CAND QL_INST_CAND0_TRSBR_31 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_31_padClk));

	CAND QL_INST_CAND0_TRSBR_32 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_32_padClk));

	CAND QL_INST_CAND0_TRSBR_33 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_33_padClk));

	CAND QL_INST_CAND1_TRSBR_29 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBR_30 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_30_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBR_31 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_31_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBR_32 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_32_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_29 (.CLKIN(nx36058z1_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx36058z1_CAND2_TRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_30 (.CLKIN(nx36058z1_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx36058z1_CAND2_TRSBR_30_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_31 (.CLKIN(nx36058z1_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx36058z1_CAND2_TRSBR_31_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_32 (.CLKIN(nx36058z1_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx36058z1_CAND2_TRSBR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBR_29 (.CLKIN(nx52746z1_SQMUX_TRSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx52746z1_CAND3_TRSBR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBR_30 (.CLKIN(nx52746z1_SQMUX_TRSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx52746z1_CAND3_TRSBR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBR_31 (.CLKIN(nx52746z1_SQMUX_TRSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx52746z1_CAND3_TRSBR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBR_32 (.CLKIN(nx52746z1_SQMUX_TRSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx52746z1_CAND3_TRSBR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSTL_0 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_0_padClk));

	CANDEN QL_INST_CAND0_BLSTL_1 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_1_padClk));

	CANDEN QL_INST_CAND0_BLSTL_3 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_3_padClk));

	CANDEN QL_INST_CAND0_BLSTL_4 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_4_padClk));

	CANDEN QL_INST_CAND0_BLSTL_5 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_5_padClk));

	CANDEN QL_INST_CAND0_BLSTL_6 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_6_padClk));

	CANDEN QL_INST_CAND0_BLSTL_7 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_7_padClk));

	CANDEN QL_INST_CAND0_BLSTL_8 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_8_padClk));

	CANDEN QL_INST_CAND1_BLSTL_1 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_3 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_4 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_5 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_6 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_7 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_8 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_1 (.CLKIN(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSTL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_3 (.CLKIN(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSTL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_5 (.CLKIN(nx9707z1_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTL_6 (.CLKIN(CLK_int_3__SQMUX_BLSTL3_padClk),.SEN(VCC),.IZ(CLK_int_3__CAND3_BLSTL_6_padClk));

	CAND QL_INST_CAND4_BLSTL_5 (.CLKIN(nx4939z1_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND4_BLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTL_6 (.CLKIN(nx4939z1_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND4_BLSTL_6_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTL_7 (.CLKIN(nx4939z1_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND4_BLSTL_7_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTL_8 (.CLKIN(nx4939z1_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND4_BLSTL_8_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_1 (.CLKIN(NET_29_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(NET_29_CAND5_BLSTL_1_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_7 (.CLKIN(NET_29_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(NET_29_CAND5_BLSTL_7_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_8 (.CLKIN(NET_29_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(NET_29_CAND5_BLSTL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSTR_9 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_9_padClk));

	CANDEN QL_INST_CAND0_BLSTR_10 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_10_padClk));

	CANDEN QL_INST_CAND0_BLSTR_11 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_11_padClk));

	CANDEN QL_INST_CAND0_BLSTR_12 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_12_padClk));

	CANDEN QL_INST_CAND0_BLSTR_13 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_13_padClk));

	CANDEN QL_INST_CAND0_BLSTR_14 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_14_padClk));

	CANDEN QL_INST_CAND0_BLSTR_15 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_15_padClk));

	CANDEN QL_INST_CAND0_BLSTR_16 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_16_padClk));

	CANDEN QL_INST_CAND1_BLSTR_9 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_10 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_11 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_12 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_13 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_14 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_15 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_16 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_9 (.CLKIN(nx19726z1_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx19726z1_CAND2_BLSTR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_10 (.CLKIN(nx19726z1_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx19726z1_CAND2_BLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_11 (.CLKIN(nx19726z1_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx19726z1_CAND2_BLSTR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_12 (.CLKIN(nx19726z1_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx19726z1_CAND2_BLSTR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_13 (.CLKIN(nx19726z1_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx19726z1_CAND2_BLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_14 (.CLKIN(nx19726z1_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx19726z1_CAND2_BLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_10 (.CLKIN(NET_17_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_17_CAND3_BLSTR_10_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_11 (.CLKIN(NET_17_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_17_CAND3_BLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_12 (.CLKIN(NET_17_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_17_CAND3_BLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_13 (.CLKIN(NET_17_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_17_CAND3_BLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_14 (.CLKIN(NET_17_SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_17_CAND3_BLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_9 (.CLKIN(NET_28_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_28_CAND4_BLSTR_9_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_10 (.CLKIN(NET_28_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_28_CAND4_BLSTR_10_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_11 (.CLKIN(NET_28_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_28_CAND4_BLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_13 (.CLKIN(NET_28_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_28_CAND4_BLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_14 (.CLKIN(NET_28_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_28_CAND4_BLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_10 (.CLKIN(NET_18_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_18_CAND5_BLSTR_10_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_11 (.CLKIN(NET_18_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_18_CAND5_BLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_12 (.CLKIN(NET_18_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_18_CAND5_BLSTR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSBL_1 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_1_padClk));

	CANDEN QL_INST_CAND0_BLSBL_2 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_2_padClk));

	CANDEN QL_INST_CAND0_BLSBL_3 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_3_padClk));

	CANDEN QL_INST_CAND0_BLSBL_4 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_4_padClk));

	CANDEN QL_INST_CAND0_BLSBL_5 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_5_padClk));

	CANDEN QL_INST_CAND0_BLSBL_6 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_6_padClk));

	CANDEN QL_INST_CAND0_BLSBL_7 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_7_padClk));

	CANDEN QL_INST_CAND0_BLSBL_8 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_8_padClk));

	CANDEN QL_INST_CAND1_BLSBL_1 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_2 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_3 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_4 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_5 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_6 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_7 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_8 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_1 (.CLKIN(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSBL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_2 (.CLKIN(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSBL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_3 (.CLKIN(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSBL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_5 (.CLKIN(nx9707z1_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx9707z1_CAND2_BLSBL_5_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBL_7 (.CLKIN(nx60831z1_SQMUX_BLSBL3_tpGCLKBUF),.SEN(VCC),.IZ(nx60831z1_CAND3_BLSBL_7_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBL_8 (.CLKIN(nx60831z1_SQMUX_BLSBL3_tpGCLKBUF),.SEN(VCC),.IZ(nx60831z1_CAND3_BLSBL_8_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBL_3 (.CLKIN(nx22245z1_SQMUX_BLSBL4_tpGCLKBUF),.SEN(VCC),.IZ(nx22245z1_CAND4_BLSBL_3_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBL_4 (.CLKIN(nx22245z1_SQMUX_BLSBL4_tpGCLKBUF),.SEN(VCC),.IZ(nx22245z1_CAND4_BLSBL_4_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBL_5 (.CLKIN(nx22245z1_SQMUX_BLSBL4_tpGCLKBUF),.SEN(VCC),.IZ(nx22245z1_CAND4_BLSBL_5_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBL_6 (.CLKIN(nx22245z1_SQMUX_BLSBL4_tpGCLKBUF),.SEN(VCC),.IZ(nx22245z1_CAND4_BLSBL_6_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBL_7 (.CLKIN(nx22245z1_SQMUX_BLSBL4_tpGCLKBUF),.SEN(VCC),.IZ(nx22245z1_CAND4_BLSBL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSBR_9 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_9_padClk));

	CANDEN QL_INST_CAND0_BLSBR_10 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_10_padClk));

	CANDEN QL_INST_CAND0_BLSBR_11 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_11_padClk));

	CANDEN QL_INST_CAND0_BLSBR_13 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_13_padClk));

	CANDEN QL_INST_CAND0_BLSBR_14 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_14_padClk));

	CANDEN QL_INST_CAND0_BLSBR_15 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_15_padClk));

	CANDEN QL_INST_CAND0_BLSBR_16 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_16_padClk));

	CANDEN QL_INST_CAND1_BLSBR_9 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_10 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_11 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_13 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_14 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_15 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_16 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_13 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_14 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_15 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_16 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_16_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_11 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_11_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_12 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_12_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_13 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_13_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_14 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_15 (.CLKIN(NET_43_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(NET_43_CAND3_BLSBR_15_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBR_12 (.CLKIN(NET_44_SQMUX_BLSBR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_44_CAND4_BLSBR_12_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBR_13 (.CLKIN(NET_44_SQMUX_BLSBR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_44_CAND4_BLSBR_13_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBR_14 (.CLKIN(NET_44_SQMUX_BLSBR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_44_CAND4_BLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBR_15 (.CLKIN(NET_44_SQMUX_BLSBR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_44_CAND4_BLSBR_15_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSBR_10 (.CLKIN(NET_32_SQMUX_BLSBR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_32_CAND5_BLSBR_10_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSBR_11 (.CLKIN(NET_32_SQMUX_BLSBR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_32_CAND5_BLSBR_11_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSBR_12 (.CLKIN(NET_32_SQMUX_BLSBR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_32_CAND5_BLSBR_12_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSBR_13 (.CLKIN(NET_32_SQMUX_BLSBR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_32_CAND5_BLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSTL_17 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_17_padClk));

	CANDEN QL_INST_CAND0_BRSTL_18 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_18_padClk));

	CANDEN QL_INST_CAND0_BRSTL_19 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_19_padClk));

	CANDEN QL_INST_CAND0_BRSTL_20 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_20_padClk));

	CANDEN QL_INST_CAND0_BRSTL_21 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_21_padClk));

	CANDEN QL_INST_CAND0_BRSTL_22 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_22_padClk));

	CANDEN QL_INST_CAND1_BRSTL_17 (.CLKIN(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTL_18 (.CLKIN(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTL_18_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTL_19 (.CLKIN(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTL_20 (.CLKIN(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTL_21 (.CLKIN(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTL_22 (.CLKIN(not_RESET_0_SQMUX_BRSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTL_22_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_18 (.CLKIN(NET_83_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_83_CAND2_BRSTL_18_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_19 (.CLKIN(NET_83_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_83_CAND2_BRSTL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_20 (.CLKIN(NET_83_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_83_CAND2_BRSTL_20_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTL_17 (.CLKIN(NET_125_SQMUX_BRSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_125_CAND3_BRSTL_17_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTL_17 (.CLKIN(NET_110_SQMUX_BRSTL4_tpGCLKBUF),.SEN(VCC),.IZ(NET_110_CAND4_BRSTL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSTR_28 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_28_padClk));

	CANDEN QL_INST_CAND0_BRSTR_29 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_29_padClk));

	CANDEN QL_INST_CAND0_BRSTR_30 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_30_padClk));

	CANDEN QL_INST_CAND0_BRSTR_31 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_31_padClk));

	CANDEN QL_INST_CAND0_BRSTR_32 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_32_padClk));

	CANDEN QL_INST_CAND0_BRSTR_33 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_33_padClk));

	CANDEN QL_INST_CAND1_BRSTR_28 (.CLKIN(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTR_29 (.CLKIN(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTR_30 (.CLKIN(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTR_31 (.CLKIN(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTR_32 (.CLKIN(not_RESET_0_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSTR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_30 (.CLKIN(nx2520z1_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSTR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_31 (.CLKIN(nx2520z1_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSTR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_32 (.CLKIN(nx2520z1_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSTR_32_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTR_30 (.CLKIN(nx57881z1_SQMUX_BRSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx57881z1_CAND3_BRSTR_30_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTR_31 (.CLKIN(nx57881z1_SQMUX_BRSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx57881z1_CAND3_BRSTR_31_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTR_32 (.CLKIN(nx57881z1_SQMUX_BRSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx57881z1_CAND3_BRSTR_32_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTR_29 (.CLKIN(nx30923z1_SQMUX_BRSTR4_tpGCLKBUF),.SEN(VCC),.IZ(nx30923z1_CAND4_BRSTR_29_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTR_30 (.CLKIN(nx30923z1_SQMUX_BRSTR4_tpGCLKBUF),.SEN(VCC),.IZ(nx30923z1_CAND4_BRSTR_30_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTR_31 (.CLKIN(nx30923z1_SQMUX_BRSTR4_tpGCLKBUF),.SEN(VCC),.IZ(nx30923z1_CAND4_BRSTR_31_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTR_32 (.CLKIN(nx30923z1_SQMUX_BRSTR4_tpGCLKBUF),.SEN(VCC),.IZ(nx30923z1_CAND4_BRSTR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSBL_17 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_17_padClk));

	CANDEN QL_INST_CAND0_BRSBL_18 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_18_padClk));

	CANDEN QL_INST_CAND0_BRSBL_19 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_19_padClk));

	CANDEN QL_INST_CAND0_BRSBL_23 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_23_padClk));

	CANDEN QL_INST_CAND0_BRSBL_24 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_24_padClk));

	CANDEN QL_INST_CAND1_BRSBL_17 (.CLKIN(not_RESET_0_SQMUX_BRSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBL_18 (.CLKIN(not_RESET_0_SQMUX_BRSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBL_18_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBL_23 (.CLKIN(not_RESET_0_SQMUX_BRSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBL_23_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBL_24 (.CLKIN(not_RESET_0_SQMUX_BRSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBL_24_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBL_17 (.CLKIN(nx14650z1_SQMUX_BRSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx14650z1_CAND2_BRSBL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBL_18 (.CLKIN(nx14650z1_SQMUX_BRSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx14650z1_CAND2_BRSBL_18_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSBR_25 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_25_padClk));

	CANDEN QL_INST_CAND0_BRSBR_26 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_26_padClk));

	CANDEN QL_INST_CAND0_BRSBR_27 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_27_padClk));

	CANDEN QL_INST_CAND0_BRSBR_28 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_28_padClk));

	CANDEN QL_INST_CAND0_BRSBR_29 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_29_padClk));

	CANDEN QL_INST_CAND0_BRSBR_30 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_30_padClk));

	CANDEN QL_INST_CAND0_BRSBR_31 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_31_padClk));

	CANDEN QL_INST_CAND0_BRSBR_32 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_32_padClk));

	CANDEN QL_INST_CAND1_BRSBR_25 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_26 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_27 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_28 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_29 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_30 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_31 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_32 (.CLKIN(not_RESET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BRSBR_32_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_30 (.CLKIN(nx2520z1_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSBR_30_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_31 (.CLKIN(nx2520z1_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSBR_31_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_32 (.CLKIN(nx2520z1_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx2520z1_CAND2_BRSBR_32_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_29 (.CLKIN(nx25788z1_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z1_CAND3_BRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_30 (.CLKIN(nx25788z1_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z1_CAND3_BRSBR_30_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_31 (.CLKIN(nx25788z1_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z1_CAND3_BRSBR_31_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_32 (.CLKIN(nx25788z1_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z1_CAND3_BRSBR_32_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBR_28 (.CLKIN(nx53672z1_SQMUX_BRSBR4_tpGCLKBUF),.SEN(VCC),.IZ(nx53672z1_CAND4_BRSBR_28_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBR_29 (.CLKIN(nx53672z1_SQMUX_BRSBR4_tpGCLKBUF),.SEN(VCC),.IZ(nx53672z1_CAND4_BRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBR_25 (.CLKIN(nx30664z1_SQMUX_BRSBR5_tpGCLKBUF),.SEN(VCC),.IZ(nx30664z1_CAND5_BRSBR_25_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBR_26 (.CLKIN(nx30664z1_SQMUX_BRSBR5_tpGCLKBUF),.SEN(VCC),.IZ(nx30664z1_CAND5_BRSBR_26_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBR_27 (.CLKIN(nx30664z1_SQMUX_BRSBR5_tpGCLKBUF),.SEN(VCC),.IZ(nx30664z1_CAND5_BRSBR_27_tpGCLKBUF));

	qlIBUF QL_INST_A2F_T_3_2 (.IN_IBUF(m0_oper0_rdata[31]),.OUT_IBUF(m0_oper0_rdata_int[31]));

	qlIBUF QL_INST_A2F_T_3_3 (.IN_IBUF(m0_oper0_rdata[30]),.OUT_IBUF(m0_oper0_rdata_int[30]));

	qlIBUF QL_INST_A2F_T_3_4 (.IN_IBUF(m0_oper0_rdata[29]),.OUT_IBUF(m0_oper0_rdata_int[29]));

	qlIBUF QL_INST_A2F_T_3_5 (.IN_IBUF(m0_oper0_rdata[28]),.OUT_IBUF(m0_oper0_rdata_int[28]));

	qlOBUF QL_INST_F2A_T_4_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTL_4_padClk),.OUT_OBUF(m0_oper0_wclk));

	qlOBUF QL_INST_F2A_T_4_2 (.IN_OBUF(m0_oper0_wmode_dup_0[1]),.OUT_OBUF(m0_oper0_wmode[1]));

	qlOBUF QL_INST_F2A_T_4_3 (.IN_OBUF(m0_oper0_wmode_dup_0[0]),.OUT_OBUF(m0_oper0_wmode[0]));

	qlOBUF QL_INST_F2A_T_4_4 (.IN_OBUF(m0_oper0_wdata_dup_0[31]),.OUT_OBUF(m0_oper0_wdata[31]));

	qlOBUF QL_INST_F2A_T_4_5 (.IN_OBUF(m0_oper0_wdata_dup_0[30]),.OUT_OBUF(m0_oper0_wdata[30]));

	qlOBUF QL_INST_F2A_T_4_6 (.IN_OBUF(m0_oper0_wdata_dup_0[29]),.OUT_OBUF(m0_oper0_wdata[29]));

	qlOBUF QL_INST_F2A_T_4_7 (.IN_OBUF(m0_oper0_wdata_dup_0[28]),.OUT_OBUF(m0_oper0_wdata[28]));

	qlOBUF QL_INST_F2A_T_4_8 (.IN_OBUF(m0_oper0_wdata_dup_0[27]),.OUT_OBUF(m0_oper0_wdata[27]));

	qlOBUF QL_INST_F2A_T_4_9 (.IN_OBUF(m0_oper0_wdata_dup_0[26]),.OUT_OBUF(m0_oper0_wdata[26]));

	qlOBUF QL_INST_F2A_T_4_10 (.IN_OBUF(m0_oper0_wdata_dup_0[25]),.OUT_OBUF(m0_oper0_wdata[25]));

	qlOBUF QL_INST_F2A_T_4_11 (.IN_OBUF(m0_oper0_wdata_dup_0[24]),.OUT_OBUF(m0_oper0_wdata[24]));

	qlOBUF QL_INST_F2A_T_4_12 (.IN_OBUF(m0_oper0_wdata_dup_0[23]),.OUT_OBUF(m0_oper0_wdata[23]));

	qlOBUF QL_INST_F2A_T_4_13 (.IN_OBUF(m0_oper0_wdata_dup_0[22]),.OUT_OBUF(m0_oper0_wdata[22]));

	qlOBUF QL_INST_F2A_T_4_14 (.IN_OBUF(m0_oper0_wdata_dup_0[21]),.OUT_OBUF(m0_oper0_wdata[21]));

	qlOBUF QL_INST_F2A_T_4_15 (.IN_OBUF(m0_oper0_wdata_dup_0[20]),.OUT_OBUF(m0_oper0_wdata[20]));

	qlOBUF QL_INST_F2A_T_4_16 (.IN_OBUF(m0_oper0_wdata_dup_0[19]),.OUT_OBUF(m0_oper0_wdata[19]));

	qlOBUF QL_INST_F2A_T_4_17 (.IN_OBUF(m0_oper0_wdata_dup_0[18]),.OUT_OBUF(m0_oper0_wdata[18]));

	qlIBUF QL_INST_A2F_T_4_0 (.IN_IBUF(m0_oper0_rdata[27]),.OUT_IBUF(m0_oper0_rdata_int[27]));

	qlIBUF QL_INST_A2F_T_4_1 (.IN_IBUF(m0_oper0_rdata[26]),.OUT_IBUF(m0_oper0_rdata_int[26]));

	qlIBUF QL_INST_A2F_T_4_2 (.IN_IBUF(m0_oper0_rdata[25]),.OUT_IBUF(m0_oper0_rdata_int[25]));

	qlIBUF QL_INST_A2F_T_4_3 (.IN_IBUF(m0_oper0_rdata[24]),.OUT_IBUF(m0_oper0_rdata_int[24]));

	qlIBUF QL_INST_A2F_T_4_4 (.IN_IBUF(m0_oper0_rdata[23]),.OUT_IBUF(m0_oper0_rdata_int[23]));

	qlIBUF QL_INST_A2F_T_4_5 (.IN_IBUF(m0_oper0_rdata[22]),.OUT_IBUF(m0_oper0_rdata_int[22]));

	qlIBUF QL_INST_A2F_T_4_6 (.IN_IBUF(m0_oper0_rdata[21]),.OUT_IBUF(m0_oper0_rdata_int[21]));

	qlIBUF QL_INST_A2F_T_4_7 (.IN_IBUF(m0_oper0_rdata[20]),.OUT_IBUF(m0_oper0_rdata_int[20]));

	qlOBUF QL_INST_F2A_T_5_0 (.IN_OBUF(m0_oper0_wdata_dup_0[17]),.OUT_OBUF(m0_oper0_wdata[17]));

	qlOBUF QL_INST_F2A_T_5_1 (.IN_OBUF(m0_oper0_wdata_dup_0[16]),.OUT_OBUF(m0_oper0_wdata[16]));

	qlOBUF QL_INST_F2A_T_5_2 (.IN_OBUF(m0_oper0_wdata_dup_0[15]),.OUT_OBUF(m0_oper0_wdata[15]));

	qlOBUF QL_INST_F2A_T_5_3 (.IN_OBUF(m0_oper0_wdata_dup_0[14]),.OUT_OBUF(m0_oper0_wdata[14]));

	qlOBUF QL_INST_F2A_T_5_4 (.IN_OBUF(m0_oper0_wdata_dup_0[13]),.OUT_OBUF(m0_oper0_wdata[13]));

	qlOBUF QL_INST_F2A_T_5_5 (.IN_OBUF(m0_oper0_wdata_dup_0[12]),.OUT_OBUF(m0_oper0_wdata[12]));

	qlOBUF QL_INST_F2A_T_5_6 (.IN_OBUF(m0_oper0_wdata_dup_0[11]),.OUT_OBUF(m0_oper0_wdata[11]));

	qlOBUF QL_INST_F2A_T_5_7 (.IN_OBUF(m0_oper0_wdata_dup_0[10]),.OUT_OBUF(m0_oper0_wdata[10]));

	qlOBUF QL_INST_F2A_T_5_8 (.IN_OBUF(m0_oper0_wdata_dup_0[9]),.OUT_OBUF(m0_oper0_wdata[9]));

	qlOBUF QL_INST_F2A_T_5_9 (.IN_OBUF(m0_oper0_wdata_dup_0[8]),.OUT_OBUF(m0_oper0_wdata[8]));

	qlOBUF QL_INST_F2A_T_5_10 (.IN_OBUF(m0_oper0_wdata_dup_0[7]),.OUT_OBUF(m0_oper0_wdata[7]));

	qlOBUF QL_INST_F2A_T_5_11 (.IN_OBUF(m0_oper0_wdata_dup_0[6]),.OUT_OBUF(m0_oper0_wdata[6]));

	qlIBUF QL_INST_A2F_T_5_0 (.IN_IBUF(m0_oper0_rdata[19]),.OUT_IBUF(m0_oper0_rdata_int[19]));

	qlIBUF QL_INST_A2F_T_5_1 (.IN_IBUF(m0_oper0_rdata[18]),.OUT_IBUF(m0_oper0_rdata_int[18]));

	qlIBUF QL_INST_A2F_T_5_2 (.IN_IBUF(m0_oper0_rdata[17]),.OUT_IBUF(m0_oper0_rdata_int[17]));

	qlIBUF QL_INST_A2F_T_5_3 (.IN_IBUF(m0_oper0_rdata[16]),.OUT_IBUF(m0_oper0_rdata_int[16]));

	qlIBUF QL_INST_A2F_T_5_4 (.IN_IBUF(m0_oper0_rdata[15]),.OUT_IBUF(m0_oper0_rdata_int[15]));

	qlIBUF QL_INST_A2F_T_5_5 (.IN_IBUF(m0_oper0_rdata[14]),.OUT_IBUF(m0_oper0_rdata_int[14]));

	qlOBUF QL_INST_F2A_T_6_0 (.IN_OBUF(m0_oper0_wdata_dup_0[5]),.OUT_OBUF(m0_oper0_wdata[5]));

	qlOBUF QL_INST_F2A_T_6_1 (.IN_OBUF(m0_oper0_wdata_dup_0[4]),.OUT_OBUF(m0_oper0_wdata[4]));

	qlOBUF QL_INST_F2A_T_6_2 (.IN_OBUF(m0_oper0_wdata_dup_0[3]),.OUT_OBUF(m0_oper0_wdata[3]));

	qlOBUF QL_INST_F2A_T_6_3 (.IN_OBUF(m0_oper0_wdata_dup_0[2]),.OUT_OBUF(m0_oper0_wdata[2]));

	qlOBUF QL_INST_F2A_T_6_4 (.IN_OBUF(m0_oper0_wdata_dup_0[1]),.OUT_OBUF(m0_oper0_wdata[1]));

	qlOBUF QL_INST_F2A_T_6_5 (.IN_OBUF(m0_oper0_wdata_dup_0[0]),.OUT_OBUF(m0_oper0_wdata[0]));

	qlOBUF QL_INST_F2A_T_6_7 (.IN_OBUF(m0_oper0_waddr_dup_0[11]),.OUT_OBUF(m0_oper0_waddr[11]));

	qlOBUF QL_INST_F2A_T_6_8 (.IN_OBUF(m0_oper0_waddr_dup_0[10]),.OUT_OBUF(m0_oper0_waddr[10]));

	qlOBUF QL_INST_F2A_T_6_9 (.IN_OBUF(m0_oper0_waddr_dup_0[9]),.OUT_OBUF(m0_oper0_waddr[9]));

	qlOBUF QL_INST_F2A_T_6_10 (.IN_OBUF(m0_oper0_waddr_dup_0[8]),.OUT_OBUF(m0_oper0_waddr[8]));

	qlOBUF QL_INST_F2A_T_6_11 (.IN_OBUF(m0_oper0_waddr_dup_0[7]),.OUT_OBUF(m0_oper0_waddr[7]));

	qlOBUF QL_INST_F2A_T_6_12 (.IN_OBUF(m0_oper0_waddr_dup_0[6]),.OUT_OBUF(m0_oper0_waddr[6]));

	qlOBUF QL_INST_F2A_T_6_13 (.IN_OBUF(m0_oper0_waddr_dup_0[5]),.OUT_OBUF(m0_oper0_waddr[5]));

	qlOBUF QL_INST_F2A_T_6_14 (.IN_OBUF(m0_oper0_waddr_dup_0[4]),.OUT_OBUF(m0_oper0_waddr[4]));

	qlOBUF QL_INST_F2A_T_6_15 (.IN_OBUF(m0_oper0_waddr_dup_0[3]),.OUT_OBUF(m0_oper0_waddr[3]));

	qlOBUF QL_INST_F2A_T_6_16 (.IN_OBUF(m0_oper0_waddr_dup_0[2]),.OUT_OBUF(m0_oper0_waddr[2]));

	qlOBUF QL_INST_F2A_T_6_17 (.IN_OBUF(m0_oper0_waddr_dup_0[1]),.OUT_OBUF(m0_oper0_waddr[1]));

	DBUF QL_INST_F2Adef_T_6_1 (.IN_DBUF(GND),.OUT_DBUF(m1_oper1_powerdn));

	qlIBUF QL_INST_A2F_T_6_0 (.IN_IBUF(m0_oper0_rdata[13]),.OUT_IBUF(m0_oper0_rdata_int[13]));

	qlIBUF QL_INST_A2F_T_6_1 (.IN_IBUF(m0_oper0_rdata[12]),.OUT_IBUF(m0_oper0_rdata_int[12]));

	qlIBUF QL_INST_A2F_T_6_2 (.IN_IBUF(m0_oper0_rdata[11]),.OUT_IBUF(m0_oper0_rdata_int[11]));

	qlIBUF QL_INST_A2F_T_6_3 (.IN_IBUF(m0_oper0_rdata[10]),.OUT_IBUF(m0_oper0_rdata_int[10]));

	qlIBUF QL_INST_A2F_T_6_4 (.IN_IBUF(m0_oper0_rdata[9]),.OUT_IBUF(m0_oper0_rdata_int[9]));

	qlIBUF QL_INST_A2F_T_6_5 (.IN_IBUF(m0_oper0_rdata[8]),.OUT_IBUF(m0_oper0_rdata_int[8]));

	qlIBUF QL_INST_A2F_T_6_6 (.IN_IBUF(m0_oper0_rdata[7]),.OUT_IBUF(m0_oper0_rdata_int[7]));

	qlIBUF QL_INST_A2F_T_6_7 (.IN_IBUF(m0_oper0_rdata[6]),.OUT_IBUF(m0_oper0_rdata_int[6]));

	qlOBUF QL_INST_F2A_T_7_0 (.IN_OBUF(m0_oper0_waddr_dup_0[0]),.OUT_OBUF(m0_oper0_waddr[0]));

	qlOBUF QL_INST_F2A_T_7_1 (.IN_OBUF(m0_oper0_we_dup_0),.OUT_OBUF(m0_oper0_we));

	qlOBUF QL_INST_F2A_T_7_2 (.IN_OBUF(m0_oper0_wdsel_dup_0),.OUT_OBUF(m0_oper0_wdsel));

	qlOBUF QL_INST_F2A_T_7_3 (.IN_OBUF(m0_oper0_rmode_dup_0[1]),.OUT_OBUF(m0_oper0_rmode[1]));

	qlOBUF QL_INST_F2A_T_7_4 (.IN_OBUF(m0_oper0_rmode_dup_0[0]),.OUT_OBUF(m0_oper0_rmode[0]));

	qlOBUF QL_INST_F2A_T_7_5 (.IN_OBUF(m0_oper0_raddr_dup_0[11]),.OUT_OBUF(m0_oper0_raddr[11]));

	qlOBUF QL_INST_F2A_T_7_6 (.IN_OBUF(m0_oper0_raddr_dup_0[10]),.OUT_OBUF(m0_oper0_raddr[10]));

	qlOBUF QL_INST_F2A_T_7_7 (.IN_OBUF(m0_oper0_raddr_dup_0[9]),.OUT_OBUF(m0_oper0_raddr[9]));

	qlOBUF QL_INST_F2A_T_7_8 (.IN_OBUF(m0_oper0_raddr_dup_0[8]),.OUT_OBUF(m0_oper0_raddr[8]));

	qlOBUF QL_INST_F2A_T_7_9 (.IN_OBUF(m0_oper0_raddr_dup_0[7]),.OUT_OBUF(m0_oper0_raddr[7]));

	qlOBUF QL_INST_F2A_T_7_10 (.IN_OBUF(m0_oper0_raddr_dup_0[6]),.OUT_OBUF(m0_oper0_raddr[6]));

	qlOBUF QL_INST_F2A_T_7_11 (.IN_OBUF(m0_oper0_raddr_dup_0[5]),.OUT_OBUF(m0_oper0_raddr[5]));

	qlIBUF QL_INST_A2F_T_7_0 (.IN_IBUF(m0_oper0_rdata[5]),.OUT_IBUF(m0_oper0_rdata_int[5]));

	qlIBUF QL_INST_A2F_T_7_1 (.IN_IBUF(m0_oper0_rdata[4]),.OUT_IBUF(m0_oper0_rdata_int[4]));

	qlIBUF QL_INST_A2F_T_7_2 (.IN_IBUF(m0_oper0_rdata[3]),.OUT_IBUF(m0_oper0_rdata_int[3]));

	qlIBUF QL_INST_A2F_T_7_3 (.IN_IBUF(m0_oper0_rdata[2]),.OUT_IBUF(m0_oper0_rdata_int[2]));

	qlIBUF QL_INST_A2F_T_7_4 (.IN_IBUF(m0_oper0_rdata[1]),.OUT_IBUF(m0_oper0_rdata_int[1]));

	qlIBUF QL_INST_A2F_T_7_5 (.IN_IBUF(m0_oper0_rdata[0]),.OUT_IBUF(m0_oper0_rdata_int[0]));

	qlOBUF QL_INST_F2A_T_8_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTL_8_padClk),.OUT_OBUF(m0_oper0_rclk));

	qlOBUF QL_INST_F2A_T_8_1 (.IN_OBUF(m0_oper0_raddr_dup_0[4]),.OUT_OBUF(m0_oper0_raddr[4]));

	qlOBUF QL_INST_F2A_T_8_2 (.IN_OBUF(m0_oper0_raddr_dup_0[3]),.OUT_OBUF(m0_oper0_raddr[3]));

	qlOBUF QL_INST_F2A_T_8_3 (.IN_OBUF(m0_oper0_raddr_dup_0[2]),.OUT_OBUF(m0_oper0_raddr[2]));

	qlOBUF QL_INST_F2A_T_8_4 (.IN_OBUF(m0_oper0_raddr_dup_0[1]),.OUT_OBUF(m0_oper0_raddr[1]));

	qlOBUF QL_INST_F2A_T_8_5 (.IN_OBUF(m0_oper0_raddr_dup_0[0]),.OUT_OBUF(m0_oper0_raddr[0]));

	qlOBUF QL_INST_F2A_T_8_7 (.IN_OBUF(m0_m0_osel_dup_0),.OUT_OBUF(m0_m0_osel));

	qlOBUF QL_INST_F2A_T_8_8 (.IN_OBUF(m0_m0_clken_dup_0),.OUT_OBUF(m0_m0_clken));

	qlOBUF QL_INST_F2A_T_8_9 (.IN_OBUF(m0_m0_outsel_dup_0[5]),.OUT_OBUF(m0_m0_outsel[5]));

	qlOBUF QL_INST_F2A_T_8_10 (.IN_OBUF(m0_m0_outsel_dup_0[4]),.OUT_OBUF(m0_m0_outsel[4]));

	qlOBUF QL_INST_F2A_T_8_11 (.IN_OBUF(m0_m0_outsel_dup_0[3]),.OUT_OBUF(m0_m0_outsel[3]));

	qlOBUF QL_INST_F2A_T_8_12 (.IN_OBUF(m0_m0_outsel_dup_0[2]),.OUT_OBUF(m0_m0_outsel[2]));

	qlOBUF QL_INST_F2A_T_8_13 (.IN_OBUF(m0_m0_outsel_dup_0[1]),.OUT_OBUF(m0_m0_outsel[1]));

	qlOBUF QL_INST_F2A_T_8_14 (.IN_OBUF(m0_m0_outsel_dup_0[0]),.OUT_OBUF(m0_m0_outsel[0]));

	qlOBUF QL_INST_F2A_T_8_15 (.IN_OBUF(m0_m0_sat_dup_0),.OUT_OBUF(m0_m0_sat));

	qlOBUF QL_INST_F2A_T_8_16 (.IN_OBUF(m0_m0_rnd_dup_0),.OUT_OBUF(m0_m0_rnd));

	qlOBUF QL_INST_F2A_T_8_17 (.IN_OBUF(m0_m0_clr_dup_0),.OUT_OBUF(m0_m0_clr));

	qlIBUF QL_INST_A2F_T_8_4 (.IN_IBUF(m0_m0_dataout[31]),.OUT_IBUF(m0_m0_dataout_int[31]));

	qlIBUF QL_INST_A2F_T_8_5 (.IN_IBUF(m0_m0_dataout[30]),.OUT_IBUF(m0_m0_dataout_int[30]));

	qlIBUF QL_INST_A2F_T_8_6 (.IN_IBUF(m0_m0_dataout[29]),.OUT_IBUF(m0_m0_dataout_int[29]));

	qlIBUF QL_INST_A2F_T_8_7 (.IN_IBUF(m0_m0_dataout[28]),.OUT_IBUF(m0_m0_dataout_int[28]));

	qlOBUF QL_INST_F2A_T_9_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTR_9_padClk),.OUT_OBUF(m0_m0_clk));

	qlOBUF QL_INST_F2A_T_9_1 (.IN_OBUF(m0_oper0_rdata_int[31]),.OUT_OBUF(m0_m0_oper_in[31]));

	qlOBUF QL_INST_F2A_T_9_2 (.IN_OBUF(m0_oper0_rdata_int[30]),.OUT_OBUF(m0_m0_oper_in[30]));

	qlOBUF QL_INST_F2A_T_9_3 (.IN_OBUF(m0_oper0_rdata_int[29]),.OUT_OBUF(m0_m0_oper_in[29]));

	qlOBUF QL_INST_F2A_T_9_4 (.IN_OBUF(m0_oper0_rdata_int[28]),.OUT_OBUF(m0_m0_oper_in[28]));

	qlOBUF QL_INST_F2A_T_9_5 (.IN_OBUF(m0_oper0_rdata_int[27]),.OUT_OBUF(m0_m0_oper_in[27]));

	qlOBUF QL_INST_F2A_T_9_6 (.IN_OBUF(m0_oper0_rdata_int[26]),.OUT_OBUF(m0_m0_oper_in[26]));

	qlOBUF QL_INST_F2A_T_9_7 (.IN_OBUF(m0_oper0_rdata_int[25]),.OUT_OBUF(m0_m0_oper_in[25]));

	qlOBUF QL_INST_F2A_T_9_8 (.IN_OBUF(m0_oper0_rdata_int[24]),.OUT_OBUF(m0_m0_oper_in[24]));

	qlOBUF QL_INST_F2A_T_9_9 (.IN_OBUF(m0_oper0_rdata_int[23]),.OUT_OBUF(m0_m0_oper_in[23]));

	qlOBUF QL_INST_F2A_T_9_10 (.IN_OBUF(m0_oper0_rdata_int[22]),.OUT_OBUF(m0_m0_oper_in[22]));

	qlOBUF QL_INST_F2A_T_9_11 (.IN_OBUF(m0_oper0_rdata_int[21]),.OUT_OBUF(m0_m0_oper_in[21]));

	qlIBUF QL_INST_A2F_T_9_0 (.IN_IBUF(m0_m0_dataout[27]),.OUT_IBUF(m0_m0_dataout_int[27]));

	qlIBUF QL_INST_A2F_T_9_1 (.IN_IBUF(m0_m0_dataout[26]),.OUT_IBUF(m0_m0_dataout_int[26]));

	qlIBUF QL_INST_A2F_T_9_2 (.IN_IBUF(m0_m0_dataout[25]),.OUT_IBUF(m0_m0_dataout_int[25]));

	qlIBUF QL_INST_A2F_T_9_3 (.IN_IBUF(m0_m0_dataout[24]),.OUT_IBUF(m0_m0_dataout_int[24]));

	qlIBUF QL_INST_A2F_T_9_4 (.IN_IBUF(m0_m0_dataout[23]),.OUT_IBUF(m0_m0_dataout_int[23]));

	qlIBUF QL_INST_A2F_T_9_5 (.IN_IBUF(m0_m0_dataout[22]),.OUT_IBUF(m0_m0_dataout_int[22]));

	qlOBUF QL_INST_F2A_T_10_0 (.IN_OBUF(m0_oper0_rdata_int[20]),.OUT_OBUF(m0_m0_oper_in[20]));

	qlOBUF QL_INST_F2A_T_10_1 (.IN_OBUF(m0_oper0_rdata_int[19]),.OUT_OBUF(m0_m0_oper_in[19]));

	qlOBUF QL_INST_F2A_T_10_2 (.IN_OBUF(m0_oper0_rdata_int[18]),.OUT_OBUF(m0_m0_oper_in[18]));

	qlOBUF QL_INST_F2A_T_10_3 (.IN_OBUF(m0_oper0_rdata_int[17]),.OUT_OBUF(m0_m0_oper_in[17]));

	qlOBUF QL_INST_F2A_T_10_4 (.IN_OBUF(m0_oper0_rdata_int[16]),.OUT_OBUF(m0_m0_oper_in[16]));

	qlOBUF QL_INST_F2A_T_10_5 (.IN_OBUF(m0_oper0_rdata_int[15]),.OUT_OBUF(m0_m0_oper_in[15]));

	qlOBUF QL_INST_F2A_T_10_6 (.IN_OBUF(m0_oper0_rdata_int[14]),.OUT_OBUF(m0_m0_oper_in[14]));

	qlOBUF QL_INST_F2A_T_10_7 (.IN_OBUF(m0_oper0_rdata_int[13]),.OUT_OBUF(m0_m0_oper_in[13]));

	qlOBUF QL_INST_F2A_T_10_8 (.IN_OBUF(m0_oper0_rdata_int[12]),.OUT_OBUF(m0_m0_oper_in[12]));

	qlOBUF QL_INST_F2A_T_10_9 (.IN_OBUF(m0_oper0_rdata_int[11]),.OUT_OBUF(m0_m0_oper_in[11]));

	qlOBUF QL_INST_F2A_T_10_10 (.IN_OBUF(m0_oper0_rdata_int[10]),.OUT_OBUF(m0_m0_oper_in[10]));

	qlOBUF QL_INST_F2A_T_10_11 (.IN_OBUF(m0_oper0_rdata_int[9]),.OUT_OBUF(m0_m0_oper_in[9]));

	qlOBUF QL_INST_F2A_T_10_12 (.IN_OBUF(m0_oper0_rdata_int[8]),.OUT_OBUF(m0_m0_oper_in[8]));

	qlOBUF QL_INST_F2A_T_10_13 (.IN_OBUF(m0_oper0_rdata_int[7]),.OUT_OBUF(m0_m0_oper_in[7]));

	qlOBUF QL_INST_F2A_T_10_14 (.IN_OBUF(m0_oper0_rdata_int[6]),.OUT_OBUF(m0_m0_oper_in[6]));

	qlOBUF QL_INST_F2A_T_10_15 (.IN_OBUF(m0_oper0_rdata_int[5]),.OUT_OBUF(m0_m0_oper_in[5]));

	qlOBUF QL_INST_F2A_T_10_16 (.IN_OBUF(m0_oper0_rdata_int[4]),.OUT_OBUF(m0_m0_oper_in[4]));

	qlOBUF QL_INST_F2A_T_10_17 (.IN_OBUF(m0_oper0_rdata_int[3]),.OUT_OBUF(m0_m0_oper_in[3]));

	qlIBUF QL_INST_A2F_T_10_0 (.IN_IBUF(m0_m0_dataout[21]),.OUT_IBUF(m0_m0_dataout_int[21]));

	qlIBUF QL_INST_A2F_T_10_1 (.IN_IBUF(m0_m0_dataout[20]),.OUT_IBUF(m0_m0_dataout_int[20]));

	qlIBUF QL_INST_A2F_T_10_2 (.IN_IBUF(m0_m0_dataout[19]),.OUT_IBUF(m0_m0_dataout_int[19]));

	qlIBUF QL_INST_A2F_T_10_3 (.IN_IBUF(m0_m0_dataout[18]),.OUT_IBUF(m0_m0_dataout_int[18]));

	qlIBUF QL_INST_A2F_T_10_4 (.IN_IBUF(m0_m0_dataout[17]),.OUT_IBUF(m0_m0_dataout_int[17]));

	qlIBUF QL_INST_A2F_T_10_5 (.IN_IBUF(m0_m0_dataout[16]),.OUT_IBUF(m0_m0_dataout_int[16]));

	qlIBUF QL_INST_A2F_T_10_6 (.IN_IBUF(m0_m0_dataout[15]),.OUT_IBUF(m0_m0_dataout_int[15]));

	qlIBUF QL_INST_A2F_T_10_7 (.IN_IBUF(m0_m0_dataout[14]),.OUT_IBUF(m0_m0_dataout_int[14]));

	qlOBUF QL_INST_F2A_T_11_0 (.IN_OBUF(m0_oper0_rdata_int[2]),.OUT_OBUF(m0_m0_oper_in[2]));

	qlOBUF QL_INST_F2A_T_11_1 (.IN_OBUF(m0_oper0_rdata_int[1]),.OUT_OBUF(m0_m0_oper_in[1]));

	qlOBUF QL_INST_F2A_T_11_2 (.IN_OBUF(m0_oper0_rdata_int[0]),.OUT_OBUF(m0_m0_oper_in[0]));

	qlOBUF QL_INST_F2A_T_11_3 (.IN_OBUF(m0_m0_csel_dup_0),.OUT_OBUF(m0_m0_csel));

	qlOBUF QL_INST_F2A_T_11_4 (.IN_OBUF(m0_coef_rdata_int[31]),.OUT_OBUF(m0_m0_coef_in[31]));

	qlOBUF QL_INST_F2A_T_11_5 (.IN_OBUF(m0_coef_rdata_int[30]),.OUT_OBUF(m0_m0_coef_in[30]));

	qlOBUF QL_INST_F2A_T_11_6 (.IN_OBUF(m0_coef_rdata_int[29]),.OUT_OBUF(m0_m0_coef_in[29]));

	qlOBUF QL_INST_F2A_T_11_7 (.IN_OBUF(m0_coef_rdata_int[28]),.OUT_OBUF(m0_m0_coef_in[28]));

	qlOBUF QL_INST_F2A_T_11_8 (.IN_OBUF(m0_coef_rdata_int[27]),.OUT_OBUF(m0_m0_coef_in[27]));

	qlOBUF QL_INST_F2A_T_11_9 (.IN_OBUF(m0_coef_rdata_int[26]),.OUT_OBUF(m0_m0_coef_in[26]));

	qlOBUF QL_INST_F2A_T_11_10 (.IN_OBUF(m0_coef_rdata_int[25]),.OUT_OBUF(m0_m0_coef_in[25]));

	qlOBUF QL_INST_F2A_T_11_11 (.IN_OBUF(m0_coef_rdata_int[24]),.OUT_OBUF(m0_m0_coef_in[24]));

	qlIBUF QL_INST_A2F_T_11_0 (.IN_IBUF(m0_m0_dataout[13]),.OUT_IBUF(m0_m0_dataout_int[13]));

	qlIBUF QL_INST_A2F_T_11_1 (.IN_IBUF(m0_m0_dataout[12]),.OUT_IBUF(m0_m0_dataout_int[12]));

	qlIBUF QL_INST_A2F_T_11_2 (.IN_IBUF(m0_m0_dataout[11]),.OUT_IBUF(m0_m0_dataout_int[11]));

	qlIBUF QL_INST_A2F_T_11_3 (.IN_IBUF(m0_m0_dataout[10]),.OUT_IBUF(m0_m0_dataout_int[10]));

	qlIBUF QL_INST_A2F_T_11_4 (.IN_IBUF(m0_m0_dataout[9]),.OUT_IBUF(m0_m0_dataout_int[9]));

	qlIBUF QL_INST_A2F_T_11_5 (.IN_IBUF(m0_m0_dataout[8]),.OUT_IBUF(m0_m0_dataout_int[8]));

	qlOBUF QL_INST_F2A_T_12_0 (.IN_OBUF(m0_coef_rdata_int[23]),.OUT_OBUF(m0_m0_coef_in[23]));

	qlOBUF QL_INST_F2A_T_12_1 (.IN_OBUF(m0_coef_rdata_int[22]),.OUT_OBUF(m0_m0_coef_in[22]));

	qlOBUF QL_INST_F2A_T_12_2 (.IN_OBUF(m0_coef_rdata_int[21]),.OUT_OBUF(m0_m0_coef_in[21]));

	qlOBUF QL_INST_F2A_T_12_3 (.IN_OBUF(m0_coef_rdata_int[20]),.OUT_OBUF(m0_m0_coef_in[20]));

	qlOBUF QL_INST_F2A_T_12_4 (.IN_OBUF(m0_coef_rdata_int[19]),.OUT_OBUF(m0_m0_coef_in[19]));

	qlOBUF QL_INST_F2A_T_12_5 (.IN_OBUF(m0_coef_rdata_int[18]),.OUT_OBUF(m0_m0_coef_in[18]));

	qlOBUF QL_INST_F2A_T_12_6 (.IN_OBUF(m0_coef_rdata_int[17]),.OUT_OBUF(m0_m0_coef_in[17]));

	qlOBUF QL_INST_F2A_T_12_7 (.IN_OBUF(m0_coef_rdata_int[16]),.OUT_OBUF(m0_m0_coef_in[16]));

	qlOBUF QL_INST_F2A_T_12_8 (.IN_OBUF(m0_coef_rdata_int[15]),.OUT_OBUF(m0_m0_coef_in[15]));

	qlOBUF QL_INST_F2A_T_12_9 (.IN_OBUF(m0_coef_rdata_int[14]),.OUT_OBUF(m0_m0_coef_in[14]));

	qlOBUF QL_INST_F2A_T_12_10 (.IN_OBUF(m0_coef_rdata_int[13]),.OUT_OBUF(m0_m0_coef_in[13]));

	qlOBUF QL_INST_F2A_T_12_11 (.IN_OBUF(m0_coef_rdata_int[12]),.OUT_OBUF(m0_m0_coef_in[12]));

	qlOBUF QL_INST_F2A_T_12_12 (.IN_OBUF(m0_coef_rdata_int[11]),.OUT_OBUF(m0_m0_coef_in[11]));

	qlOBUF QL_INST_F2A_T_12_13 (.IN_OBUF(m0_coef_rdata_int[10]),.OUT_OBUF(m0_m0_coef_in[10]));

	qlOBUF QL_INST_F2A_T_12_14 (.IN_OBUF(m0_coef_rdata_int[9]),.OUT_OBUF(m0_m0_coef_in[9]));

	qlOBUF QL_INST_F2A_T_12_15 (.IN_OBUF(m0_coef_rdata_int[8]),.OUT_OBUF(m0_m0_coef_in[8]));

	qlOBUF QL_INST_F2A_T_12_16 (.IN_OBUF(m0_coef_rdata_int[7]),.OUT_OBUF(m0_m0_coef_in[7]));

	qlOBUF QL_INST_F2A_T_12_17 (.IN_OBUF(m0_coef_rdata_int[6]),.OUT_OBUF(m0_m0_coef_in[6]));

	qlIBUF QL_INST_A2F_T_12_0 (.IN_IBUF(m0_m0_dataout[7]),.OUT_IBUF(m0_m0_dataout_int[7]));

	qlIBUF QL_INST_A2F_T_12_1 (.IN_IBUF(m0_m0_dataout[6]),.OUT_IBUF(m0_m0_dataout_int[6]));

	qlIBUF QL_INST_A2F_T_12_2 (.IN_IBUF(m0_m0_dataout[5]),.OUT_IBUF(m0_m0_dataout_int[5]));

	qlIBUF QL_INST_A2F_T_12_3 (.IN_IBUF(m0_m0_dataout[4]),.OUT_IBUF(m0_m0_dataout_int[4]));

	qlIBUF QL_INST_A2F_T_12_4 (.IN_IBUF(m0_m0_dataout[3]),.OUT_IBUF(m0_m0_dataout_int[3]));

	qlIBUF QL_INST_A2F_T_12_5 (.IN_IBUF(m0_m0_dataout[2]),.OUT_IBUF(m0_m0_dataout_int[2]));

	qlIBUF QL_INST_A2F_T_12_6 (.IN_IBUF(m0_m0_dataout[1]),.OUT_IBUF(m0_m0_dataout_int[1]));

	qlIBUF QL_INST_A2F_T_12_7 (.IN_IBUF(m0_m0_dataout[0]),.OUT_IBUF(m0_m0_dataout_int[0]));

	qlOBUF QL_INST_F2A_T_13_0 (.IN_OBUF(m0_coef_rdata_int[5]),.OUT_OBUF(m0_m0_coef_in[5]));

	qlOBUF QL_INST_F2A_T_13_1 (.IN_OBUF(m0_coef_rdata_int[4]),.OUT_OBUF(m0_m0_coef_in[4]));

	qlOBUF QL_INST_F2A_T_13_2 (.IN_OBUF(m0_coef_rdata_int[3]),.OUT_OBUF(m0_m0_coef_in[3]));

	qlOBUF QL_INST_F2A_T_13_3 (.IN_OBUF(m0_coef_rdata_int[2]),.OUT_OBUF(m0_m0_coef_in[2]));

	qlOBUF QL_INST_F2A_T_13_4 (.IN_OBUF(m0_coef_rdata_int[1]),.OUT_OBUF(m0_m0_coef_in[1]));

	qlOBUF QL_INST_F2A_T_13_5 (.IN_OBUF(m0_coef_rdata_int[0]),.OUT_OBUF(m0_m0_coef_in[0]));

	qlOBUF QL_INST_F2A_T_13_6 (.IN_OBUF(m0_m0_mode_dup_0[1]),.OUT_OBUF(m0_m0_mode[1]));

	qlOBUF QL_INST_F2A_T_13_7 (.IN_OBUF(m0_m0_mode_dup_0[0]),.OUT_OBUF(m0_m0_mode[0]));

	qlOBUF QL_INST_F2A_T_13_8 (.IN_OBUF(m0_m0_tc_dup_0),.OUT_OBUF(m0_m0_tc));

	qlOBUF QL_INST_F2A_T_13_9 (.IN_OBUF(m0_m0_reset_dup_0),.OUT_OBUF(m0_m0_reset));

	qlOBUF QL_INST_F2A_T_13_10 (.IN_OBUF(m0_coef_wdata_dup_0[31]),.OUT_OBUF(m0_coef_wdata[31]));

	qlOBUF QL_INST_F2A_T_13_11 (.IN_OBUF(m0_coef_wdata_dup_0[30]),.OUT_OBUF(m0_coef_wdata[30]));

	DBUF QL_INST_F2Adef_T_13_0 (.IN_DBUF(GND),.OUT_DBUF(m1_coef_powerdn));

	qlIBUF QL_INST_A2F_T_13_2 (.IN_IBUF(m0_coef_rdata[31]),.OUT_IBUF(m0_coef_rdata_int[31]));

	qlIBUF QL_INST_A2F_T_13_3 (.IN_IBUF(m0_coef_rdata[30]),.OUT_IBUF(m0_coef_rdata_int[30]));

	qlIBUF QL_INST_A2F_T_13_4 (.IN_IBUF(m0_coef_rdata[29]),.OUT_IBUF(m0_coef_rdata_int[29]));

	qlIBUF QL_INST_A2F_T_13_5 (.IN_IBUF(m0_coef_rdata[28]),.OUT_IBUF(m0_coef_rdata_int[28]));

	qlOBUF QL_INST_F2A_T_14_0 (.IN_OBUF(m0_coef_wdata_dup_0[29]),.OUT_OBUF(m0_coef_wdata[29]));

	qlOBUF QL_INST_F2A_T_14_1 (.IN_OBUF(m0_coef_wdata_dup_0[28]),.OUT_OBUF(m0_coef_wdata[28]));

	qlOBUF QL_INST_F2A_T_14_2 (.IN_OBUF(m0_coef_wdata_dup_0[27]),.OUT_OBUF(m0_coef_wdata[27]));

	qlOBUF QL_INST_F2A_T_14_3 (.IN_OBUF(m0_coef_wdata_dup_0[26]),.OUT_OBUF(m0_coef_wdata[26]));

	qlOBUF QL_INST_F2A_T_14_4 (.IN_OBUF(m0_coef_wdata_dup_0[25]),.OUT_OBUF(m0_coef_wdata[25]));

	qlOBUF QL_INST_F2A_T_14_5 (.IN_OBUF(m0_coef_wdata_dup_0[24]),.OUT_OBUF(m0_coef_wdata[24]));

	qlOBUF QL_INST_F2A_T_14_6 (.IN_OBUF(m0_coef_wdata_dup_0[23]),.OUT_OBUF(m0_coef_wdata[23]));

	qlOBUF QL_INST_F2A_T_14_7 (.IN_OBUF(m0_coef_wdata_dup_0[22]),.OUT_OBUF(m0_coef_wdata[22]));

	qlOBUF QL_INST_F2A_T_14_8 (.IN_OBUF(m0_coef_wdata_dup_0[21]),.OUT_OBUF(m0_coef_wdata[21]));

	qlOBUF QL_INST_F2A_T_14_9 (.IN_OBUF(m0_coef_wdata_dup_0[20]),.OUT_OBUF(m0_coef_wdata[20]));

	qlOBUF QL_INST_F2A_T_14_10 (.IN_OBUF(m0_coef_wdata_dup_0[19]),.OUT_OBUF(m0_coef_wdata[19]));

	qlOBUF QL_INST_F2A_T_14_11 (.IN_OBUF(m0_coef_wdata_dup_0[18]),.OUT_OBUF(m0_coef_wdata[18]));

	qlOBUF QL_INST_F2A_T_14_12 (.IN_OBUF(m0_coef_wdata_dup_0[17]),.OUT_OBUF(m0_coef_wdata[17]));

	qlOBUF QL_INST_F2A_T_14_13 (.IN_OBUF(m0_coef_wdata_dup_0[16]),.OUT_OBUF(m0_coef_wdata[16]));

	qlOBUF QL_INST_F2A_T_14_14 (.IN_OBUF(m0_coef_wdata_dup_0[15]),.OUT_OBUF(m0_coef_wdata[15]));

	qlOBUF QL_INST_F2A_T_14_15 (.IN_OBUF(m0_coef_wdata_dup_0[14]),.OUT_OBUF(m0_coef_wdata[14]));

	qlOBUF QL_INST_F2A_T_14_16 (.IN_OBUF(m0_coef_wdata_dup_0[13]),.OUT_OBUF(m0_coef_wdata[13]));

	qlOBUF QL_INST_F2A_T_14_17 (.IN_OBUF(m0_coef_wdata_dup_0[12]),.OUT_OBUF(m0_coef_wdata[12]));

	qlIBUF QL_INST_A2F_T_14_0 (.IN_IBUF(m0_coef_rdata[27]),.OUT_IBUF(m0_coef_rdata_int[27]));

	qlIBUF QL_INST_A2F_T_14_1 (.IN_IBUF(m0_coef_rdata[26]),.OUT_IBUF(m0_coef_rdata_int[26]));

	qlIBUF QL_INST_A2F_T_14_2 (.IN_IBUF(m0_coef_rdata[25]),.OUT_IBUF(m0_coef_rdata_int[25]));

	qlIBUF QL_INST_A2F_T_14_3 (.IN_IBUF(m0_coef_rdata[24]),.OUT_IBUF(m0_coef_rdata_int[24]));

	qlIBUF QL_INST_A2F_T_14_4 (.IN_IBUF(m0_coef_rdata[23]),.OUT_IBUF(m0_coef_rdata_int[23]));

	qlIBUF QL_INST_A2F_T_14_5 (.IN_IBUF(m0_coef_rdata[22]),.OUT_IBUF(m0_coef_rdata_int[22]));

	qlIBUF QL_INST_A2F_T_14_6 (.IN_IBUF(m0_coef_rdata[21]),.OUT_IBUF(m0_coef_rdata_int[21]));

	qlIBUF QL_INST_A2F_T_14_7 (.IN_IBUF(m0_coef_rdata[20]),.OUT_IBUF(m0_coef_rdata_int[20]));

	qlOBUF QL_INST_F2A_T_15_0 (.IN_OBUF(m0_coef_wdata_dup_0[11]),.OUT_OBUF(m0_coef_wdata[11]));

	qlOBUF QL_INST_F2A_T_15_1 (.IN_OBUF(m0_coef_wdata_dup_0[10]),.OUT_OBUF(m0_coef_wdata[10]));

	qlOBUF QL_INST_F2A_T_15_2 (.IN_OBUF(m0_coef_wdata_dup_0[9]),.OUT_OBUF(m0_coef_wdata[9]));

	qlOBUF QL_INST_F2A_T_15_3 (.IN_OBUF(m0_coef_wdata_dup_0[8]),.OUT_OBUF(m0_coef_wdata[8]));

	qlOBUF QL_INST_F2A_T_15_4 (.IN_OBUF(m0_coef_wdata_dup_0[7]),.OUT_OBUF(m0_coef_wdata[7]));

	qlOBUF QL_INST_F2A_T_15_5 (.IN_OBUF(m0_coef_wdata_dup_0[6]),.OUT_OBUF(m0_coef_wdata[6]));

	qlOBUF QL_INST_F2A_T_15_6 (.IN_OBUF(m0_coef_wdata_dup_0[5]),.OUT_OBUF(m0_coef_wdata[5]));

	qlOBUF QL_INST_F2A_T_15_7 (.IN_OBUF(m0_coef_wdata_dup_0[4]),.OUT_OBUF(m0_coef_wdata[4]));

	qlOBUF QL_INST_F2A_T_15_8 (.IN_OBUF(m0_coef_wdata_dup_0[3]),.OUT_OBUF(m0_coef_wdata[3]));

	qlOBUF QL_INST_F2A_T_15_9 (.IN_OBUF(m0_coef_wdata_dup_0[2]),.OUT_OBUF(m0_coef_wdata[2]));

	qlOBUF QL_INST_F2A_T_15_10 (.IN_OBUF(m0_coef_wdata_dup_0[1]),.OUT_OBUF(m0_coef_wdata[1]));

	qlOBUF QL_INST_F2A_T_15_11 (.IN_OBUF(m0_coef_wdata_dup_0[0]),.OUT_OBUF(m0_coef_wdata[0]));

	qlIBUF QL_INST_A2F_T_15_0 (.IN_IBUF(m0_coef_rdata[19]),.OUT_IBUF(m0_coef_rdata_int[19]));

	qlIBUF QL_INST_A2F_T_15_1 (.IN_IBUF(m0_coef_rdata[18]),.OUT_IBUF(m0_coef_rdata_int[18]));

	qlIBUF QL_INST_A2F_T_15_2 (.IN_IBUF(m0_coef_rdata[17]),.OUT_IBUF(m0_coef_rdata_int[17]));

	qlIBUF QL_INST_A2F_T_15_3 (.IN_IBUF(m0_coef_rdata[16]),.OUT_IBUF(m0_coef_rdata_int[16]));

	qlIBUF QL_INST_A2F_T_15_4 (.IN_IBUF(m0_coef_rdata[15]),.OUT_IBUF(m0_coef_rdata_int[15]));

	qlIBUF QL_INST_A2F_T_15_5 (.IN_IBUF(m0_coef_rdata[14]),.OUT_IBUF(m0_coef_rdata_int[14]));

	qlOBUF QL_INST_F2A_T_16_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTR_16_padClk),.OUT_OBUF(m0_coef_wclk));

	qlOBUF QL_INST_F2A_T_16_1 (.IN_OBUF(m0_coef_waddr_dup_0[11]),.OUT_OBUF(m0_coef_waddr[11]));

	qlOBUF QL_INST_F2A_T_16_2 (.IN_OBUF(m0_coef_waddr_dup_0[10]),.OUT_OBUF(m0_coef_waddr[10]));

	qlOBUF QL_INST_F2A_T_16_3 (.IN_OBUF(m0_coef_waddr_dup_0[9]),.OUT_OBUF(m0_coef_waddr[9]));

	qlOBUF QL_INST_F2A_T_16_4 (.IN_OBUF(m0_coef_waddr_dup_0[8]),.OUT_OBUF(m0_coef_waddr[8]));

	qlOBUF QL_INST_F2A_T_16_5 (.IN_OBUF(m0_coef_waddr_dup_0[7]),.OUT_OBUF(m0_coef_waddr[7]));

	qlOBUF QL_INST_F2A_T_16_6 (.IN_OBUF(m0_coef_waddr_dup_0[6]),.OUT_OBUF(m0_coef_waddr[6]));

	qlOBUF QL_INST_F2A_T_16_7 (.IN_OBUF(m0_coef_waddr_dup_0[5]),.OUT_OBUF(m0_coef_waddr[5]));

	qlOBUF QL_INST_F2A_T_16_8 (.IN_OBUF(m0_coef_waddr_dup_0[4]),.OUT_OBUF(m0_coef_waddr[4]));

	qlOBUF QL_INST_F2A_T_16_9 (.IN_OBUF(m0_coef_waddr_dup_0[3]),.OUT_OBUF(m0_coef_waddr[3]));

	qlOBUF QL_INST_F2A_T_16_10 (.IN_OBUF(m0_coef_waddr_dup_0[2]),.OUT_OBUF(m0_coef_waddr[2]));

	qlOBUF QL_INST_F2A_T_16_11 (.IN_OBUF(m0_coef_waddr_dup_0[1]),.OUT_OBUF(m0_coef_waddr[1]));

	qlOBUF QL_INST_F2A_T_16_12 (.IN_OBUF(m0_coef_waddr_dup_0[0]),.OUT_OBUF(m0_coef_waddr[0]));

	qlOBUF QL_INST_F2A_T_16_13 (.IN_OBUF(m0_coef_we_dup_0),.OUT_OBUF(m0_coef_we));

	qlOBUF QL_INST_F2A_T_16_17 (.IN_OBUF(m0_coef_wdsel_dup_0),.OUT_OBUF(m0_coef_wdsel));

	qlIBUF QL_INST_A2F_T_16_0 (.IN_IBUF(m0_coef_rdata[13]),.OUT_IBUF(m0_coef_rdata_int[13]));

	qlIBUF QL_INST_A2F_T_16_1 (.IN_IBUF(m0_coef_rdata[12]),.OUT_IBUF(m0_coef_rdata_int[12]));

	qlIBUF QL_INST_A2F_T_16_2 (.IN_IBUF(m0_coef_rdata[11]),.OUT_IBUF(m0_coef_rdata_int[11]));

	qlIBUF QL_INST_A2F_T_16_3 (.IN_IBUF(m0_coef_rdata[10]),.OUT_IBUF(m0_coef_rdata_int[10]));

	qlIBUF QL_INST_A2F_T_16_4 (.IN_IBUF(m0_coef_rdata[9]),.OUT_IBUF(m0_coef_rdata_int[9]));

	qlIBUF QL_INST_A2F_T_16_5 (.IN_IBUF(m0_coef_rdata[8]),.OUT_IBUF(m0_coef_rdata_int[8]));

	qlIBUF QL_INST_A2F_T_16_6 (.IN_IBUF(m0_coef_rdata[7]),.OUT_IBUF(m0_coef_rdata_int[7]));

	qlIBUF QL_INST_A2F_T_16_7 (.IN_IBUF(m0_coef_rdata[6]),.OUT_IBUF(m0_coef_rdata_int[6]));

	qlOBUF QL_INST_F2A_T_17_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTL_17_padClk),.OUT_OBUF(m0_coef_rclk));

	qlOBUF QL_INST_F2A_T_17_1 (.IN_OBUF(m0_coef_rmode_dup_0[1]),.OUT_OBUF(m0_coef_rmode[1]));

	qlOBUF QL_INST_F2A_T_17_2 (.IN_OBUF(m0_coef_rmode_dup_0[0]),.OUT_OBUF(m0_coef_rmode[0]));

	qlOBUF QL_INST_F2A_T_17_3 (.IN_OBUF(m0_coef_raddr_dup_0[11]),.OUT_OBUF(m0_coef_raddr[11]));

	qlOBUF QL_INST_F2A_T_17_4 (.IN_OBUF(m0_coef_raddr_dup_0[10]),.OUT_OBUF(m0_coef_raddr[10]));

	qlOBUF QL_INST_F2A_T_17_5 (.IN_OBUF(m0_coef_raddr_dup_0[9]),.OUT_OBUF(m0_coef_raddr[9]));

	qlOBUF QL_INST_F2A_T_17_6 (.IN_OBUF(m0_coef_raddr_dup_0[8]),.OUT_OBUF(m0_coef_raddr[8]));

	qlOBUF QL_INST_F2A_T_17_7 (.IN_OBUF(m0_coef_raddr_dup_0[7]),.OUT_OBUF(m0_coef_raddr[7]));

	qlOBUF QL_INST_F2A_T_17_8 (.IN_OBUF(m0_coef_raddr_dup_0[6]),.OUT_OBUF(m0_coef_raddr[6]));

	qlOBUF QL_INST_F2A_T_17_9 (.IN_OBUF(m0_coef_raddr_dup_0[5]),.OUT_OBUF(m0_coef_raddr[5]));

	qlOBUF QL_INST_F2A_T_17_10 (.IN_OBUF(m0_coef_raddr_dup_0[4]),.OUT_OBUF(m0_coef_raddr[4]));

	qlOBUF QL_INST_F2A_T_17_11 (.IN_OBUF(m0_coef_raddr_dup_0[3]),.OUT_OBUF(m0_coef_raddr[3]));

	qlIBUF QL_INST_A2F_T_17_0 (.IN_IBUF(m0_coef_rdata[5]),.OUT_IBUF(m0_coef_rdata_int[5]));

	qlIBUF QL_INST_A2F_T_17_1 (.IN_IBUF(m0_coef_rdata[4]),.OUT_IBUF(m0_coef_rdata_int[4]));

	qlIBUF QL_INST_A2F_T_17_2 (.IN_IBUF(m0_coef_rdata[3]),.OUT_IBUF(m0_coef_rdata_int[3]));

	qlIBUF QL_INST_A2F_T_17_3 (.IN_IBUF(m0_coef_rdata[2]),.OUT_IBUF(m0_coef_rdata_int[2]));

	qlIBUF QL_INST_A2F_T_17_4 (.IN_IBUF(m0_coef_rdata[1]),.OUT_IBUF(m0_coef_rdata_int[1]));

	qlIBUF QL_INST_A2F_T_17_5 (.IN_IBUF(m0_coef_rdata[0]),.OUT_IBUF(m0_coef_rdata_int[0]));

	qlOBUF QL_INST_F2A_T_18_1 (.IN_OBUF(m0_coef_raddr_dup_0[2]),.OUT_OBUF(m0_coef_raddr[2]));

	qlOBUF QL_INST_F2A_T_18_2 (.IN_OBUF(m0_coef_raddr_dup_0[1]),.OUT_OBUF(m0_coef_raddr[1]));

	qlOBUF QL_INST_F2A_T_18_3 (.IN_OBUF(m0_coef_raddr_dup_0[0]),.OUT_OBUF(m0_coef_raddr[0]));

	qlOBUF QL_INST_F2A_T_18_4 (.IN_OBUF(m0_coef_wmode_dup_0[1]),.OUT_OBUF(m0_coef_wmode[1]));

	qlOBUF QL_INST_F2A_T_18_5 (.IN_OBUF(m0_coef_wmode_dup_0[0]),.OUT_OBUF(m0_coef_wmode[0]));

	qlOBUF QL_INST_F2A_T_18_8 (.IN_OBUF(m0_m1_outsel_dup_0[5]),.OUT_OBUF(m0_m1_outsel[5]));

	qlOBUF QL_INST_F2A_T_18_9 (.IN_OBUF(m0_m1_outsel_dup_0[4]),.OUT_OBUF(m0_m1_outsel[4]));

	qlOBUF QL_INST_F2A_T_18_10 (.IN_OBUF(m0_m1_outsel_dup_0[3]),.OUT_OBUF(m0_m1_outsel[3]));

	qlOBUF QL_INST_F2A_T_18_11 (.IN_OBUF(m0_m1_outsel_dup_0[2]),.OUT_OBUF(m0_m1_outsel[2]));

	qlOBUF QL_INST_F2A_T_18_12 (.IN_OBUF(m0_m1_outsel_dup_0[1]),.OUT_OBUF(m0_m1_outsel[1]));

	qlOBUF QL_INST_F2A_T_18_13 (.IN_OBUF(m0_m1_outsel_dup_0[0]),.OUT_OBUF(m0_m1_outsel[0]));

	qlOBUF QL_INST_F2A_T_18_14 (.IN_OBUF(m0_m1_sat_dup_0),.OUT_OBUF(m0_m1_sat));

	qlOBUF QL_INST_F2A_T_18_15 (.IN_OBUF(m0_m1_rnd_dup_0),.OUT_OBUF(m0_m1_rnd));

	qlOBUF QL_INST_F2A_T_18_16 (.IN_OBUF(m0_m1_clr_dup_0),.OUT_OBUF(m0_m1_clr));

	qlOBUF QL_INST_F2A_T_18_17 (.IN_OBUF(m0_m1_clken_dup_0),.OUT_OBUF(m0_m1_clken));

	qlIBUF QL_INST_A2F_T_18_0 (.IN_IBUF(m0_m1_dataout[31]),.OUT_IBUF(m0_m1_dataout_int[31]));

	qlIBUF QL_INST_A2F_T_18_1 (.IN_IBUF(m0_m1_dataout[30]),.OUT_IBUF(m0_m1_dataout_int[30]));

	qlIBUF QL_INST_A2F_T_18_2 (.IN_IBUF(m0_m1_dataout[29]),.OUT_IBUF(m0_m1_dataout_int[29]));

	qlIBUF QL_INST_A2F_T_18_3 (.IN_IBUF(m0_m1_dataout[28]),.OUT_IBUF(m0_m1_dataout_int[28]));

	qlIBUF QL_INST_A2F_T_18_4 (.IN_IBUF(m0_m1_dataout[27]),.OUT_IBUF(m0_m1_dataout_int[27]));

	qlIBUF QL_INST_A2F_T_18_5 (.IN_IBUF(m0_m1_dataout[26]),.OUT_IBUF(m0_m1_dataout_int[26]));

	qlIBUF QL_INST_A2F_T_18_6 (.IN_IBUF(m0_m1_dataout[25]),.OUT_IBUF(m0_m1_dataout_int[25]));

	qlIBUF QL_INST_A2F_T_18_7 (.IN_IBUF(m0_m1_dataout[24]),.OUT_IBUF(m0_m1_dataout_int[24]));

	qlOBUF QL_INST_F2A_T_19_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTL_19_padClk),.OUT_OBUF(m0_m1_clk));

	qlOBUF QL_INST_F2A_T_19_1 (.IN_OBUF(m0_m1_osel_dup_0),.OUT_OBUF(m0_m1_osel));

	qlOBUF QL_INST_F2A_T_19_2 (.IN_OBUF(m0_m1_tc_dup_0),.OUT_OBUF(m0_m1_tc));

	qlOBUF QL_INST_F2A_T_19_3 (.IN_OBUF(m0_m1_reset_dup_0),.OUT_OBUF(m0_m1_reset));

	qlOBUF QL_INST_F2A_T_19_4 (.IN_OBUF(m0_coef_rdata_int[31]),.OUT_OBUF(m0_m1_coef_in[31]));

	qlOBUF QL_INST_F2A_T_19_5 (.IN_OBUF(m0_coef_rdata_int[30]),.OUT_OBUF(m0_m1_coef_in[30]));

	qlOBUF QL_INST_F2A_T_19_6 (.IN_OBUF(m0_coef_rdata_int[29]),.OUT_OBUF(m0_m1_coef_in[29]));

	qlOBUF QL_INST_F2A_T_19_7 (.IN_OBUF(m0_coef_rdata_int[28]),.OUT_OBUF(m0_m1_coef_in[28]));

	qlOBUF QL_INST_F2A_T_19_8 (.IN_OBUF(m0_coef_rdata_int[27]),.OUT_OBUF(m0_m1_coef_in[27]));

	qlOBUF QL_INST_F2A_T_19_9 (.IN_OBUF(m0_coef_rdata_int[26]),.OUT_OBUF(m0_m1_coef_in[26]));

	qlOBUF QL_INST_F2A_T_19_10 (.IN_OBUF(m0_coef_rdata_int[25]),.OUT_OBUF(m0_m1_coef_in[25]));

	qlOBUF QL_INST_F2A_T_19_11 (.IN_OBUF(m0_coef_rdata_int[24]),.OUT_OBUF(m0_m1_coef_in[24]));

	qlIBUF QL_INST_A2F_T_19_0 (.IN_IBUF(m0_m1_dataout[23]),.OUT_IBUF(m0_m1_dataout_int[23]));

	qlIBUF QL_INST_A2F_T_19_1 (.IN_IBUF(m0_m1_dataout[22]),.OUT_IBUF(m0_m1_dataout_int[22]));

	qlIBUF QL_INST_A2F_T_19_2 (.IN_IBUF(m0_m1_dataout[21]),.OUT_IBUF(m0_m1_dataout_int[21]));

	qlIBUF QL_INST_A2F_T_19_3 (.IN_IBUF(m0_m1_dataout[20]),.OUT_IBUF(m0_m1_dataout_int[20]));

	qlIBUF QL_INST_A2F_T_19_4 (.IN_IBUF(m0_m1_dataout[19]),.OUT_IBUF(m0_m1_dataout_int[19]));

	qlIBUF QL_INST_A2F_T_19_5 (.IN_IBUF(m0_m1_dataout[18]),.OUT_IBUF(m0_m1_dataout_int[18]));

	qlOBUF QL_INST_F2A_T_20_0 (.IN_OBUF(m0_coef_rdata_int[23]),.OUT_OBUF(m0_m1_coef_in[23]));

	qlOBUF QL_INST_F2A_T_20_1 (.IN_OBUF(m0_coef_rdata_int[22]),.OUT_OBUF(m0_m1_coef_in[22]));

	qlOBUF QL_INST_F2A_T_20_2 (.IN_OBUF(m0_coef_rdata_int[21]),.OUT_OBUF(m0_m1_coef_in[21]));

	qlOBUF QL_INST_F2A_T_20_3 (.IN_OBUF(m0_coef_rdata_int[20]),.OUT_OBUF(m0_m1_coef_in[20]));

	qlOBUF QL_INST_F2A_T_20_4 (.IN_OBUF(m0_coef_rdata_int[19]),.OUT_OBUF(m0_m1_coef_in[19]));

	qlOBUF QL_INST_F2A_T_20_5 (.IN_OBUF(m0_coef_rdata_int[18]),.OUT_OBUF(m0_m1_coef_in[18]));

	qlOBUF QL_INST_F2A_T_20_6 (.IN_OBUF(m0_coef_rdata_int[17]),.OUT_OBUF(m0_m1_coef_in[17]));

	qlOBUF QL_INST_F2A_T_20_7 (.IN_OBUF(m0_coef_rdata_int[16]),.OUT_OBUF(m0_m1_coef_in[16]));

	qlOBUF QL_INST_F2A_T_20_8 (.IN_OBUF(m0_coef_rdata_int[15]),.OUT_OBUF(m0_m1_coef_in[15]));

	qlOBUF QL_INST_F2A_T_20_9 (.IN_OBUF(m0_coef_rdata_int[14]),.OUT_OBUF(m0_m1_coef_in[14]));

	qlOBUF QL_INST_F2A_T_20_10 (.IN_OBUF(m0_coef_rdata_int[13]),.OUT_OBUF(m0_m1_coef_in[13]));

	qlOBUF QL_INST_F2A_T_20_11 (.IN_OBUF(m0_coef_rdata_int[12]),.OUT_OBUF(m0_m1_coef_in[12]));

	qlOBUF QL_INST_F2A_T_20_12 (.IN_OBUF(m0_coef_rdata_int[11]),.OUT_OBUF(m0_m1_coef_in[11]));

	qlOBUF QL_INST_F2A_T_20_13 (.IN_OBUF(m0_coef_rdata_int[10]),.OUT_OBUF(m0_m1_coef_in[10]));

	qlOBUF QL_INST_F2A_T_20_14 (.IN_OBUF(m0_coef_rdata_int[9]),.OUT_OBUF(m0_m1_coef_in[9]));

	qlOBUF QL_INST_F2A_T_20_15 (.IN_OBUF(m0_coef_rdata_int[8]),.OUT_OBUF(m0_m1_coef_in[8]));

	qlOBUF QL_INST_F2A_T_20_16 (.IN_OBUF(m0_coef_rdata_int[7]),.OUT_OBUF(m0_m1_coef_in[7]));

	qlOBUF QL_INST_F2A_T_20_17 (.IN_OBUF(m0_coef_rdata_int[6]),.OUT_OBUF(m0_m1_coef_in[6]));

	qlIBUF QL_INST_A2F_T_20_0 (.IN_IBUF(m0_m1_dataout[17]),.OUT_IBUF(m0_m1_dataout_int[17]));

	qlIBUF QL_INST_A2F_T_20_1 (.IN_IBUF(m0_m1_dataout[16]),.OUT_IBUF(m0_m1_dataout_int[16]));

	qlIBUF QL_INST_A2F_T_20_2 (.IN_IBUF(m0_m1_dataout[15]),.OUT_IBUF(m0_m1_dataout_int[15]));

	qlIBUF QL_INST_A2F_T_20_3 (.IN_IBUF(m0_m1_dataout[14]),.OUT_IBUF(m0_m1_dataout_int[14]));

	qlIBUF QL_INST_A2F_T_20_4 (.IN_IBUF(m0_m1_dataout[13]),.OUT_IBUF(m0_m1_dataout_int[13]));

	qlIBUF QL_INST_A2F_T_20_5 (.IN_IBUF(m0_m1_dataout[12]),.OUT_IBUF(m0_m1_dataout_int[12]));

	qlIBUF QL_INST_A2F_T_20_6 (.IN_IBUF(m0_m1_dataout[11]),.OUT_IBUF(m0_m1_dataout_int[11]));

	qlOBUF QL_INST_F2A_T_21_0 (.IN_OBUF(m0_coef_rdata_int[5]),.OUT_OBUF(m0_m1_coef_in[5]));

	qlOBUF QL_INST_F2A_T_21_1 (.IN_OBUF(m0_coef_rdata_int[4]),.OUT_OBUF(m0_m1_coef_in[4]));

	qlOBUF QL_INST_F2A_T_21_2 (.IN_OBUF(m0_coef_rdata_int[3]),.OUT_OBUF(m0_m1_coef_in[3]));

	qlOBUF QL_INST_F2A_T_21_3 (.IN_OBUF(m0_coef_rdata_int[2]),.OUT_OBUF(m0_m1_coef_in[2]));

	qlOBUF QL_INST_F2A_T_21_4 (.IN_OBUF(m0_coef_rdata_int[1]),.OUT_OBUF(m0_m1_coef_in[1]));

	qlOBUF QL_INST_F2A_T_21_5 (.IN_OBUF(m0_coef_rdata_int[0]),.OUT_OBUF(m0_m1_coef_in[0]));

	qlOBUF QL_INST_F2A_T_21_6 (.IN_OBUF(m0_m1_mode_dup_0[1]),.OUT_OBUF(m0_m1_mode[1]));

	qlOBUF QL_INST_F2A_T_21_7 (.IN_OBUF(m0_m1_csel_dup_0),.OUT_OBUF(m0_m1_csel));

	qlOBUF QL_INST_F2A_T_21_8 (.IN_OBUF(m0_m1_mode_dup_0[0]),.OUT_OBUF(m0_m1_mode[0]));

	qlOBUF QL_INST_F2A_T_21_9 (.IN_OBUF(m0_oper1_rdata_int[31]),.OUT_OBUF(m0_m1_oper_in[31]));

	qlOBUF QL_INST_F2A_T_21_10 (.IN_OBUF(m0_oper1_rdata_int[30]),.OUT_OBUF(m0_m1_oper_in[30]));

	qlOBUF QL_INST_F2A_T_21_11 (.IN_OBUF(m0_oper1_rdata_int[29]),.OUT_OBUF(m0_m1_oper_in[29]));

	qlIBUF QL_INST_A2F_T_21_0 (.IN_IBUF(m0_m1_dataout[10]),.OUT_IBUF(m0_m1_dataout_int[10]));

	qlIBUF QL_INST_A2F_T_21_1 (.IN_IBUF(m0_m1_dataout[9]),.OUT_IBUF(m0_m1_dataout_int[9]));

	qlIBUF QL_INST_A2F_T_21_2 (.IN_IBUF(m0_m1_dataout[8]),.OUT_IBUF(m0_m1_dataout_int[8]));

	qlIBUF QL_INST_A2F_T_21_3 (.IN_IBUF(m0_m1_dataout[7]),.OUT_IBUF(m0_m1_dataout_int[7]));

	qlIBUF QL_INST_A2F_T_21_4 (.IN_IBUF(m0_m1_dataout[6]),.OUT_IBUF(m0_m1_dataout_int[6]));

	qlIBUF QL_INST_A2F_T_21_5 (.IN_IBUF(m0_m1_dataout[5]),.OUT_IBUF(m0_m1_dataout_int[5]));

	qlOBUF QL_INST_F2A_T_22_0 (.IN_OBUF(m0_oper1_rdata_int[28]),.OUT_OBUF(m0_m1_oper_in[28]));

	qlOBUF QL_INST_F2A_T_22_1 (.IN_OBUF(m0_oper1_rdata_int[27]),.OUT_OBUF(m0_m1_oper_in[27]));

	qlOBUF QL_INST_F2A_T_22_2 (.IN_OBUF(m0_oper1_rdata_int[26]),.OUT_OBUF(m0_m1_oper_in[26]));

	qlOBUF QL_INST_F2A_T_22_3 (.IN_OBUF(m0_oper1_rdata_int[25]),.OUT_OBUF(m0_m1_oper_in[25]));

	qlOBUF QL_INST_F2A_T_22_4 (.IN_OBUF(m0_oper1_rdata_int[24]),.OUT_OBUF(m0_m1_oper_in[24]));

	qlOBUF QL_INST_F2A_T_22_5 (.IN_OBUF(m0_oper1_rdata_int[23]),.OUT_OBUF(m0_m1_oper_in[23]));

	qlOBUF QL_INST_F2A_T_22_6 (.IN_OBUF(m0_oper1_rdata_int[22]),.OUT_OBUF(m0_m1_oper_in[22]));

	qlOBUF QL_INST_F2A_T_22_7 (.IN_OBUF(m0_oper1_rdata_int[21]),.OUT_OBUF(m0_m1_oper_in[21]));

	qlOBUF QL_INST_F2A_T_22_8 (.IN_OBUF(m0_oper1_rdata_int[20]),.OUT_OBUF(m0_m1_oper_in[20]));

	qlOBUF QL_INST_F2A_T_22_9 (.IN_OBUF(m0_oper1_rdata_int[19]),.OUT_OBUF(m0_m1_oper_in[19]));

	qlOBUF QL_INST_F2A_T_22_10 (.IN_OBUF(m0_oper1_rdata_int[18]),.OUT_OBUF(m0_m1_oper_in[18]));

	qlOBUF QL_INST_F2A_T_22_11 (.IN_OBUF(m0_oper1_rdata_int[17]),.OUT_OBUF(m0_m1_oper_in[17]));

	qlOBUF QL_INST_F2A_T_22_12 (.IN_OBUF(m0_oper1_rdata_int[16]),.OUT_OBUF(m0_m1_oper_in[16]));

	qlOBUF QL_INST_F2A_T_22_13 (.IN_OBUF(m0_oper1_rdata_int[15]),.OUT_OBUF(m0_m1_oper_in[15]));

	qlOBUF QL_INST_F2A_T_22_14 (.IN_OBUF(m0_oper1_rdata_int[14]),.OUT_OBUF(m0_m1_oper_in[14]));

	qlOBUF QL_INST_F2A_T_22_15 (.IN_OBUF(m0_oper1_rdata_int[13]),.OUT_OBUF(m0_m1_oper_in[13]));

	qlOBUF QL_INST_F2A_T_22_16 (.IN_OBUF(m0_oper1_rdata_int[12]),.OUT_OBUF(m0_m1_oper_in[12]));

	qlOBUF QL_INST_F2A_T_22_17 (.IN_OBUF(m0_oper1_rdata_int[11]),.OUT_OBUF(m0_m1_oper_in[11]));

	qlIBUF QL_INST_A2F_T_22_0 (.IN_IBUF(m0_m1_dataout[4]),.OUT_IBUF(m0_m1_dataout_int[4]));

	qlIBUF QL_INST_A2F_T_22_1 (.IN_IBUF(m0_m1_dataout[3]),.OUT_IBUF(m0_m1_dataout_int[3]));

	qlIBUF QL_INST_A2F_T_22_2 (.IN_IBUF(m0_m1_dataout[2]),.OUT_IBUF(m0_m1_dataout_int[2]));

	qlIBUF QL_INST_A2F_T_22_3 (.IN_IBUF(m0_m1_dataout[1]),.OUT_IBUF(m0_m1_dataout_int[1]));

	qlIBUF QL_INST_A2F_T_22_4 (.IN_IBUF(m0_m1_dataout[0]),.OUT_IBUF(m0_m1_dataout_int[0]));

	qlOBUF QL_INST_F2A_T_23_0 (.IN_OBUF(m0_oper1_rdata_int[10]),.OUT_OBUF(m0_m1_oper_in[10]));

	qlOBUF QL_INST_F2A_T_23_1 (.IN_OBUF(m0_oper1_rdata_int[9]),.OUT_OBUF(m0_m1_oper_in[9]));

	qlOBUF QL_INST_F2A_T_23_2 (.IN_OBUF(m0_oper1_rdata_int[8]),.OUT_OBUF(m0_m1_oper_in[8]));

	qlOBUF QL_INST_F2A_T_23_3 (.IN_OBUF(m0_oper1_rdata_int[7]),.OUT_OBUF(m0_m1_oper_in[7]));

	qlOBUF QL_INST_F2A_T_23_4 (.IN_OBUF(m0_oper1_rdata_int[6]),.OUT_OBUF(m0_m1_oper_in[6]));

	qlOBUF QL_INST_F2A_T_23_5 (.IN_OBUF(m0_oper1_rdata_int[5]),.OUT_OBUF(m0_m1_oper_in[5]));

	qlOBUF QL_INST_F2A_T_23_6 (.IN_OBUF(m0_oper1_rdata_int[4]),.OUT_OBUF(m0_m1_oper_in[4]));

	qlOBUF QL_INST_F2A_T_23_7 (.IN_OBUF(m0_oper1_rdata_int[3]),.OUT_OBUF(m0_m1_oper_in[3]));

	qlOBUF QL_INST_F2A_T_23_8 (.IN_OBUF(m0_oper1_rdata_int[2]),.OUT_OBUF(m0_m1_oper_in[2]));

	qlOBUF QL_INST_F2A_T_23_9 (.IN_OBUF(m0_oper1_rdata_int[1]),.OUT_OBUF(m0_m1_oper_in[1]));

	qlOBUF QL_INST_F2A_T_23_10 (.IN_OBUF(m0_oper1_rdata_int[0]),.OUT_OBUF(m0_m1_oper_in[0]));

	qlOBUF QL_INST_F2A_T_24_16 (.IN_OBUF(m0_oper1_wdata_dup_0[31]),.OUT_OBUF(m0_oper1_wdata[31]));

	qlOBUF QL_INST_F2A_T_24_17 (.IN_OBUF(m0_oper1_wdata_dup_0[30]),.OUT_OBUF(m0_oper1_wdata[30]));

	DBUF QL_INST_F2Adef_T_24_0 (.IN_DBUF(GND),.OUT_DBUF(m1_oper0_powerdn));

	qlOBUF QL_INST_F2A_T_25_0 (.IN_OBUF(m0_oper1_wdata_dup_0[29]),.OUT_OBUF(m0_oper1_wdata[29]));

	qlOBUF QL_INST_F2A_T_25_1 (.IN_OBUF(m0_oper1_wdata_dup_0[28]),.OUT_OBUF(m0_oper1_wdata[28]));

	qlOBUF QL_INST_F2A_T_25_2 (.IN_OBUF(m0_oper1_wdata_dup_0[27]),.OUT_OBUF(m0_oper1_wdata[27]));

	qlOBUF QL_INST_F2A_T_25_3 (.IN_OBUF(m0_oper1_wdata_dup_0[26]),.OUT_OBUF(m0_oper1_wdata[26]));

	qlOBUF QL_INST_F2A_T_25_4 (.IN_OBUF(m0_oper1_wdata_dup_0[25]),.OUT_OBUF(m0_oper1_wdata[25]));

	qlOBUF QL_INST_F2A_T_25_5 (.IN_OBUF(m0_oper1_wdata_dup_0[24]),.OUT_OBUF(m0_oper1_wdata[24]));

	qlOBUF QL_INST_F2A_T_25_6 (.IN_OBUF(m0_oper1_wdata_dup_0[23]),.OUT_OBUF(m0_oper1_wdata[23]));

	qlOBUF QL_INST_F2A_T_25_7 (.IN_OBUF(m0_oper1_wdata_dup_0[22]),.OUT_OBUF(m0_oper1_wdata[22]));

	qlOBUF QL_INST_F2A_T_25_8 (.IN_OBUF(m0_oper1_wdata_dup_0[21]),.OUT_OBUF(m0_oper1_wdata[21]));

	qlOBUF QL_INST_F2A_T_25_9 (.IN_OBUF(m0_oper1_wdata_dup_0[20]),.OUT_OBUF(m0_oper1_wdata[20]));

	qlOBUF QL_INST_F2A_T_25_10 (.IN_OBUF(m0_oper1_wdata_dup_0[19]),.OUT_OBUF(m0_oper1_wdata[19]));

	qlOBUF QL_INST_F2A_T_25_11 (.IN_OBUF(m0_oper1_wdata_dup_0[18]),.OUT_OBUF(m0_oper1_wdata[18]));

	qlIBUF QL_INST_A2F_T_25_1 (.IN_IBUF(m0_oper1_rdata[31]),.OUT_IBUF(m0_oper1_rdata_int[31]));

	qlIBUF QL_INST_A2F_T_25_2 (.IN_IBUF(m0_oper1_rdata[30]),.OUT_IBUF(m0_oper1_rdata_int[30]));

	qlIBUF QL_INST_A2F_T_25_3 (.IN_IBUF(m0_oper1_rdata[29]),.OUT_IBUF(m0_oper1_rdata_int[29]));

	qlIBUF QL_INST_A2F_T_25_4 (.IN_IBUF(m0_oper1_rdata[28]),.OUT_IBUF(m0_oper1_rdata_int[28]));

	qlIBUF QL_INST_A2F_T_25_5 (.IN_IBUF(m0_oper1_rdata[27]),.OUT_IBUF(m0_oper1_rdata_int[27]));

	qlOBUF QL_INST_F2A_T_26_0 (.IN_OBUF(m0_oper1_wdata_dup_0[17]),.OUT_OBUF(m0_oper1_wdata[17]));

	qlOBUF QL_INST_F2A_T_26_1 (.IN_OBUF(m0_oper1_wdata_dup_0[16]),.OUT_OBUF(m0_oper1_wdata[16]));

	qlOBUF QL_INST_F2A_T_26_2 (.IN_OBUF(m0_oper1_wdata_dup_0[15]),.OUT_OBUF(m0_oper1_wdata[15]));

	qlOBUF QL_INST_F2A_T_26_3 (.IN_OBUF(m0_oper1_wdata_dup_0[14]),.OUT_OBUF(m0_oper1_wdata[14]));

	qlOBUF QL_INST_F2A_T_26_4 (.IN_OBUF(m0_oper1_wdata_dup_0[13]),.OUT_OBUF(m0_oper1_wdata[13]));

	qlOBUF QL_INST_F2A_T_26_5 (.IN_OBUF(m0_oper1_wdata_dup_0[12]),.OUT_OBUF(m0_oper1_wdata[12]));

	qlOBUF QL_INST_F2A_T_26_6 (.IN_OBUF(m0_oper1_wdata_dup_0[11]),.OUT_OBUF(m0_oper1_wdata[11]));

	qlOBUF QL_INST_F2A_T_26_7 (.IN_OBUF(m0_oper1_wdata_dup_0[10]),.OUT_OBUF(m0_oper1_wdata[10]));

	qlOBUF QL_INST_F2A_T_26_8 (.IN_OBUF(m0_oper1_wdata_dup_0[9]),.OUT_OBUF(m0_oper1_wdata[9]));

	qlOBUF QL_INST_F2A_T_26_9 (.IN_OBUF(m0_oper1_wdata_dup_0[8]),.OUT_OBUF(m0_oper1_wdata[8]));

	qlOBUF QL_INST_F2A_T_26_10 (.IN_OBUF(m0_oper1_wdata_dup_0[7]),.OUT_OBUF(m0_oper1_wdata[7]));

	qlOBUF QL_INST_F2A_T_26_11 (.IN_OBUF(m0_oper1_wdata_dup_0[6]),.OUT_OBUF(m0_oper1_wdata[6]));

	qlOBUF QL_INST_F2A_T_26_12 (.IN_OBUF(m0_oper1_wdata_dup_0[5]),.OUT_OBUF(m0_oper1_wdata[5]));

	qlOBUF QL_INST_F2A_T_26_13 (.IN_OBUF(m0_oper1_wdata_dup_0[4]),.OUT_OBUF(m0_oper1_wdata[4]));

	qlOBUF QL_INST_F2A_T_26_14 (.IN_OBUF(m0_oper1_wdata_dup_0[3]),.OUT_OBUF(m0_oper1_wdata[3]));

	qlOBUF QL_INST_F2A_T_26_15 (.IN_OBUF(m0_oper1_wdata_dup_0[2]),.OUT_OBUF(m0_oper1_wdata[2]));

	qlOBUF QL_INST_F2A_T_26_16 (.IN_OBUF(m0_oper1_wdata_dup_0[1]),.OUT_OBUF(m0_oper1_wdata[1]));

	qlOBUF QL_INST_F2A_T_26_17 (.IN_OBUF(m0_oper1_wdata_dup_0[0]),.OUT_OBUF(m0_oper1_wdata[0]));

	qlIBUF QL_INST_A2F_T_26_0 (.IN_IBUF(m0_oper1_rdata[26]),.OUT_IBUF(m0_oper1_rdata_int[26]));

	qlIBUF QL_INST_A2F_T_26_1 (.IN_IBUF(m0_oper1_rdata[25]),.OUT_IBUF(m0_oper1_rdata_int[25]));

	qlIBUF QL_INST_A2F_T_26_2 (.IN_IBUF(m0_oper1_rdata[24]),.OUT_IBUF(m0_oper1_rdata_int[24]));

	qlIBUF QL_INST_A2F_T_26_3 (.IN_IBUF(m0_oper1_rdata[23]),.OUT_IBUF(m0_oper1_rdata_int[23]));

	qlIBUF QL_INST_A2F_T_26_4 (.IN_IBUF(m0_oper1_rdata[22]),.OUT_IBUF(m0_oper1_rdata_int[22]));

	qlIBUF QL_INST_A2F_T_26_5 (.IN_IBUF(m0_oper1_rdata[21]),.OUT_IBUF(m0_oper1_rdata_int[21]));

	qlIBUF QL_INST_A2F_T_26_6 (.IN_IBUF(m0_oper1_rdata[20]),.OUT_IBUF(m0_oper1_rdata_int[20]));

	qlIBUF QL_INST_A2F_T_26_7 (.IN_IBUF(m0_oper1_rdata[19]),.OUT_IBUF(m0_oper1_rdata_int[19]));

	qlOBUF QL_INST_F2A_T_27_0 (.IN_OBUF(m0_oper1_waddr_dup_0[11]),.OUT_OBUF(m0_oper1_waddr[11]));

	qlOBUF QL_INST_F2A_T_27_1 (.IN_OBUF(m0_oper1_waddr_dup_0[10]),.OUT_OBUF(m0_oper1_waddr[10]));

	qlOBUF QL_INST_F2A_T_27_2 (.IN_OBUF(m0_oper1_waddr_dup_0[9]),.OUT_OBUF(m0_oper1_waddr[9]));

	qlOBUF QL_INST_F2A_T_27_3 (.IN_OBUF(m0_oper1_waddr_dup_0[8]),.OUT_OBUF(m0_oper1_waddr[8]));

	qlOBUF QL_INST_F2A_T_27_4 (.IN_OBUF(m0_oper1_waddr_dup_0[7]),.OUT_OBUF(m0_oper1_waddr[7]));

	qlOBUF QL_INST_F2A_T_27_5 (.IN_OBUF(m0_oper1_waddr_dup_0[6]),.OUT_OBUF(m0_oper1_waddr[6]));

	qlOBUF QL_INST_F2A_T_27_6 (.IN_OBUF(m0_oper1_waddr_dup_0[5]),.OUT_OBUF(m0_oper1_waddr[5]));

	qlOBUF QL_INST_F2A_T_27_7 (.IN_OBUF(m0_oper1_waddr_dup_0[4]),.OUT_OBUF(m0_oper1_waddr[4]));

	qlOBUF QL_INST_F2A_T_27_8 (.IN_OBUF(m0_oper1_waddr_dup_0[3]),.OUT_OBUF(m0_oper1_waddr[3]));

	qlOBUF QL_INST_F2A_T_27_9 (.IN_OBUF(m0_oper1_waddr_dup_0[2]),.OUT_OBUF(m0_oper1_waddr[2]));

	qlOBUF QL_INST_F2A_T_27_10 (.IN_OBUF(m0_oper1_waddr_dup_0[1]),.OUT_OBUF(m0_oper1_waddr[1]));

	qlOBUF QL_INST_F2A_T_27_11 (.IN_OBUF(m0_oper1_waddr_dup_0[0]),.OUT_OBUF(m0_oper1_waddr[0]));

	qlIBUF QL_INST_A2F_T_27_0 (.IN_IBUF(m0_oper1_rdata[18]),.OUT_IBUF(m0_oper1_rdata_int[18]));

	qlIBUF QL_INST_A2F_T_27_1 (.IN_IBUF(m0_oper1_rdata[17]),.OUT_IBUF(m0_oper1_rdata_int[17]));

	qlIBUF QL_INST_A2F_T_27_2 (.IN_IBUF(m0_oper1_rdata[16]),.OUT_IBUF(m0_oper1_rdata_int[16]));

	qlIBUF QL_INST_A2F_T_27_3 (.IN_IBUF(m0_oper1_rdata[15]),.OUT_IBUF(m0_oper1_rdata_int[15]));

	qlIBUF QL_INST_A2F_T_27_4 (.IN_IBUF(m0_oper1_rdata[14]),.OUT_IBUF(m0_oper1_rdata_int[14]));

	qlIBUF QL_INST_A2F_T_27_5 (.IN_IBUF(m0_oper1_rdata[13]),.OUT_IBUF(m0_oper1_rdata_int[13]));

	qlOBUF QL_INST_F2A_T_28_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_28_padClk),.OUT_OBUF(m0_oper1_wclk));

	qlOBUF QL_INST_F2A_T_28_1 (.IN_OBUF(m0_oper1_wmode_dup_0[1]),.OUT_OBUF(m0_oper1_wmode[1]));

	qlOBUF QL_INST_F2A_T_28_2 (.IN_OBUF(m0_oper1_wmode_dup_0[0]),.OUT_OBUF(m0_oper1_wmode[0]));

	qlOBUF QL_INST_F2A_T_28_3 (.IN_OBUF(m0_oper1_wdsel_dup_0),.OUT_OBUF(m0_oper1_wdsel));

	qlOBUF QL_INST_F2A_T_28_4 (.IN_OBUF(m0_oper1_we_dup_0),.OUT_OBUF(m0_oper1_we));

	qlOBUF QL_INST_F2A_T_28_15 (.IN_OBUF(m0_oper1_rmode_dup_0[1]),.OUT_OBUF(m0_oper1_rmode[1]));

	qlOBUF QL_INST_F2A_T_28_16 (.IN_OBUF(m0_oper1_rmode_dup_0[0]),.OUT_OBUF(m0_oper1_rmode[0]));

	qlOBUF QL_INST_F2A_T_28_17 (.IN_OBUF(m0_oper1_raddr_dup_0[11]),.OUT_OBUF(m0_oper1_raddr[11]));

	qlIBUF QL_INST_A2F_T_28_1 (.IN_IBUF(m0_oper1_rdata[12]),.OUT_IBUF(m0_oper1_rdata_int[12]));

	qlIBUF QL_INST_A2F_T_28_2 (.IN_IBUF(m0_oper1_rdata[11]),.OUT_IBUF(m0_oper1_rdata_int[11]));

	qlIBUF QL_INST_A2F_T_28_3 (.IN_IBUF(m0_oper1_rdata[10]),.OUT_IBUF(m0_oper1_rdata_int[10]));

	qlIBUF QL_INST_A2F_T_28_4 (.IN_IBUF(m0_oper1_rdata[9]),.OUT_IBUF(m0_oper1_rdata_int[9]));

	qlIBUF QL_INST_A2F_T_28_5 (.IN_IBUF(m0_oper1_rdata[8]),.OUT_IBUF(m0_oper1_rdata_int[8]));

	qlIBUF QL_INST_A2F_T_28_6 (.IN_IBUF(m0_oper1_rdata[7]),.OUT_IBUF(m0_oper1_rdata_int[7]));

	qlIBUF QL_INST_A2F_T_28_7 (.IN_IBUF(m0_oper1_rdata[6]),.OUT_IBUF(m0_oper1_rdata_int[6]));

	qlOBUF QL_INST_F2A_T_29_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_29_padClk),.OUT_OBUF(m0_oper1_rclk));

	qlOBUF QL_INST_F2A_T_29_1 (.IN_OBUF(m0_oper1_raddr_dup_0[10]),.OUT_OBUF(m0_oper1_raddr[10]));

	qlOBUF QL_INST_F2A_T_29_2 (.IN_OBUF(m0_oper1_raddr_dup_0[9]),.OUT_OBUF(m0_oper1_raddr[9]));

	qlOBUF QL_INST_F2A_T_29_3 (.IN_OBUF(m0_oper1_raddr_dup_0[8]),.OUT_OBUF(m0_oper1_raddr[8]));

	qlOBUF QL_INST_F2A_T_29_4 (.IN_OBUF(m0_oper1_raddr_dup_0[7]),.OUT_OBUF(m0_oper1_raddr[7]));

	qlOBUF QL_INST_F2A_T_29_5 (.IN_OBUF(m0_oper1_raddr_dup_0[6]),.OUT_OBUF(m0_oper1_raddr[6]));

	qlOBUF QL_INST_F2A_T_29_6 (.IN_OBUF(m0_oper1_raddr_dup_0[5]),.OUT_OBUF(m0_oper1_raddr[5]));

	qlOBUF QL_INST_F2A_T_29_7 (.IN_OBUF(m0_oper1_raddr_dup_0[4]),.OUT_OBUF(m0_oper1_raddr[4]));

	qlOBUF QL_INST_F2A_T_29_8 (.IN_OBUF(m0_oper1_raddr_dup_0[3]),.OUT_OBUF(m0_oper1_raddr[3]));

	qlOBUF QL_INST_F2A_T_29_9 (.IN_OBUF(m0_oper1_raddr_dup_0[2]),.OUT_OBUF(m0_oper1_raddr[2]));

	qlOBUF QL_INST_F2A_T_29_10 (.IN_OBUF(m0_oper1_raddr_dup_0[1]),.OUT_OBUF(m0_oper1_raddr[1]));

	qlOBUF QL_INST_F2A_T_29_11 (.IN_OBUF(m0_oper1_raddr_dup_0[0]),.OUT_OBUF(m0_oper1_raddr[0]));

	qlIBUF QL_INST_A2F_T_29_0 (.IN_IBUF(m0_oper1_rdata[5]),.OUT_IBUF(m0_oper1_rdata_int[5]));

	qlIBUF QL_INST_A2F_T_29_1 (.IN_IBUF(m0_oper1_rdata[4]),.OUT_IBUF(m0_oper1_rdata_int[4]));

	qlIBUF QL_INST_A2F_T_29_2 (.IN_IBUF(m0_oper1_rdata[3]),.OUT_IBUF(m0_oper1_rdata_int[3]));

	qlIBUF QL_INST_A2F_T_29_3 (.IN_IBUF(m0_oper1_rdata[2]),.OUT_IBUF(m0_oper1_rdata_int[2]));

	qlIBUF QL_INST_A2F_T_29_4 (.IN_IBUF(m0_oper1_rdata[1]),.OUT_IBUF(m0_oper1_rdata_int[1]));

	qlIBUF QL_INST_A2F_T_29_5 (.IN_IBUF(m0_oper1_rdata[0]),.OUT_IBUF(m0_oper1_rdata_int[0]));

	qlOBUF QL_INST_F2A_R_3_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_33_padClk),.OUT_OBUF(tcdm_clk_p0));

	qlOBUF QL_INST_F2A_R_3_1 (.IN_OBUF(tcdm_req_p0_dup_0),.OUT_OBUF(tcdm_req_p0));

	qlOBUF QL_INST_F2A_R_3_2 (.IN_OBUF(tcdm_we_p0_dup_0),.OUT_OBUF(tcdm_we_p0));

	qlOBUF QL_INST_F2A_R_3_3 (.IN_OBUF(tcdm_be_p0_dup_0[0]),.OUT_OBUF(tcdm_be_p0[0]));

	qlOBUF QL_INST_F2A_R_3_4 (.IN_OBUF(tcdm_be_p0_dup_0[1]),.OUT_OBUF(tcdm_be_p0[1]));

	qlOBUF QL_INST_F2A_R_3_5 (.IN_OBUF(tcdm_be_p0_dup_0[2]),.OUT_OBUF(tcdm_be_p0[2]));

	qlOBUF QL_INST_F2A_R_3_6 (.IN_OBUF(tcdm_be_p0_dup_0[3]),.OUT_OBUF(tcdm_be_p0[3]));

	qlOBUF QL_INST_F2A_R_3_8 (.IN_OBUF(tcdm_addr_p0_dup_0[0]),.OUT_OBUF(tcdm_addr_p0[0]));

	qlOBUF QL_INST_F2A_R_3_9 (.IN_OBUF(tcdm_addr_p0_dup_0[1]),.OUT_OBUF(tcdm_addr_p0[1]));

	qlOBUF QL_INST_F2A_R_3_10 (.IN_OBUF(tcdm_addr_p0_dup_0[2]),.OUT_OBUF(tcdm_addr_p0[2]));

	qlOBUF QL_INST_F2A_R_3_11 (.IN_OBUF(tcdm_addr_p0_dup_0[3]),.OUT_OBUF(tcdm_addr_p0[3]));

	qlIBUF QL_INST_A2F_R_3_0 (.IN_IBUF(tcdm_rdata_p0[0]),.OUT_IBUF(tcdm_rdata_p0_int[0]));

	qlIBUF QL_INST_A2F_R_3_1 (.IN_IBUF(tcdm_rdata_p0[1]),.OUT_IBUF(tcdm_rdata_p0_int[1]));

	qlIBUF QL_INST_A2F_R_3_2 (.IN_IBUF(tcdm_rdata_p0[2]),.OUT_IBUF(tcdm_rdata_p0_int[2]));

	qlIBUF QL_INST_A2F_R_3_3 (.IN_IBUF(tcdm_rdata_p0[3]),.OUT_IBUF(tcdm_rdata_p0_int[3]));

	qlIBUF QL_INST_A2F_R_3_4 (.IN_IBUF(tcdm_valid_p0),.OUT_IBUF(tcdm_valid_p0_int));

	qlIBUF QL_INST_A2F_R_3_5 (.IN_IBUF(tcdm_gnt_p0),.OUT_IBUF(tcdm_gnt_p0_int));

	qlOBUF QL_INST_F2A_R_4_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[0]),.OUT_OBUF(tcdm_wdata_p0[0]));

	qlOBUF QL_INST_F2A_R_4_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[1]),.OUT_OBUF(tcdm_wdata_p0[1]));

	qlOBUF QL_INST_F2A_R_4_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[2]),.OUT_OBUF(tcdm_wdata_p0[2]));

	qlOBUF QL_INST_F2A_R_4_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[3]),.OUT_OBUF(tcdm_wdata_p0[3]));

	qlOBUF QL_INST_F2A_R_4_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[4]),.OUT_OBUF(tcdm_wdata_p0[4]));

	qlOBUF QL_INST_F2A_R_4_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[5]),.OUT_OBUF(tcdm_wdata_p0[5]));

	qlOBUF QL_INST_F2A_R_4_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[6]),.OUT_OBUF(tcdm_wdata_p0[6]));

	qlOBUF QL_INST_F2A_R_4_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[7]),.OUT_OBUF(tcdm_wdata_p0[7]));

	qlOBUF QL_INST_F2A_R_4_9 (.IN_OBUF(tcdm_addr_p0_dup_0[4]),.OUT_OBUF(tcdm_addr_p0[4]));

	qlOBUF QL_INST_F2A_R_4_10 (.IN_OBUF(tcdm_addr_p0_dup_0[5]),.OUT_OBUF(tcdm_addr_p0[5]));

	qlOBUF QL_INST_F2A_R_4_11 (.IN_OBUF(tcdm_addr_p0_dup_0[6]),.OUT_OBUF(tcdm_addr_p0[6]));

	qlOBUF QL_INST_F2A_R_4_12 (.IN_OBUF(tcdm_addr_p0_dup_0[7]),.OUT_OBUF(tcdm_addr_p0[7]));

	qlOBUF QL_INST_F2A_R_4_13 (.IN_OBUF(tcdm_addr_p0_dup_0[8]),.OUT_OBUF(tcdm_addr_p0[8]));

	qlOBUF QL_INST_F2A_R_4_14 (.IN_OBUF(tcdm_addr_p0_dup_0[9]),.OUT_OBUF(tcdm_addr_p0[9]));

	qlIBUF QL_INST_A2F_R_4_0 (.IN_IBUF(tcdm_rdata_p0[4]),.OUT_IBUF(tcdm_rdata_p0_int[4]));

	qlIBUF QL_INST_A2F_R_4_1 (.IN_IBUF(tcdm_rdata_p0[5]),.OUT_IBUF(tcdm_rdata_p0_int[5]));

	qlIBUF QL_INST_A2F_R_4_2 (.IN_IBUF(tcdm_rdata_p0[6]),.OUT_IBUF(tcdm_rdata_p0_int[6]));

	qlIBUF QL_INST_A2F_R_4_3 (.IN_IBUF(tcdm_rdata_p0[7]),.OUT_IBUF(tcdm_rdata_p0_int[7]));

	qlIBUF QL_INST_A2F_R_4_4 (.IN_IBUF(tcdm_rdata_p0[8]),.OUT_IBUF(tcdm_rdata_p0_int[8]));

	qlIBUF QL_INST_A2F_R_4_5 (.IN_IBUF(tcdm_rdata_p0[9]),.OUT_IBUF(tcdm_rdata_p0_int[9]));

	qlIBUF QL_INST_A2F_R_4_6 (.IN_IBUF(tcdm_rdata_p0[10]),.OUT_IBUF(tcdm_rdata_p0_int[10]));

	qlIBUF QL_INST_A2F_R_4_7 (.IN_IBUF(tcdm_rdata_p0[11]),.OUT_IBUF(tcdm_rdata_p0_int[11]));

	qlOBUF QL_INST_F2A_R_5_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[8]),.OUT_OBUF(tcdm_wdata_p0[8]));

	qlOBUF QL_INST_F2A_R_5_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[9]),.OUT_OBUF(tcdm_wdata_p0[9]));

	qlOBUF QL_INST_F2A_R_5_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[10]),.OUT_OBUF(tcdm_wdata_p0[10]));

	qlOBUF QL_INST_F2A_R_5_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[11]),.OUT_OBUF(tcdm_wdata_p0[11]));

	qlOBUF QL_INST_F2A_R_5_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[12]),.OUT_OBUF(tcdm_wdata_p0[12]));

	qlOBUF QL_INST_F2A_R_5_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[13]),.OUT_OBUF(tcdm_wdata_p0[13]));

	qlOBUF QL_INST_F2A_R_5_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[14]),.OUT_OBUF(tcdm_wdata_p0[14]));

	qlOBUF QL_INST_F2A_R_5_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[15]),.OUT_OBUF(tcdm_wdata_p0[15]));

	qlOBUF QL_INST_F2A_R_5_8 (.IN_OBUF(tcdm_addr_p0_dup_0[10]),.OUT_OBUF(tcdm_addr_p0[10]));

	qlOBUF QL_INST_F2A_R_5_9 (.IN_OBUF(tcdm_addr_p0_dup_0[11]),.OUT_OBUF(tcdm_addr_p0[11]));

	qlOBUF QL_INST_F2A_R_5_10 (.IN_OBUF(tcdm_addr_p0_dup_0[12]),.OUT_OBUF(tcdm_addr_p0[12]));

	qlOBUF QL_INST_F2A_R_5_11 (.IN_OBUF(tcdm_addr_p0_dup_0[13]),.OUT_OBUF(tcdm_addr_p0[13]));

	qlIBUF QL_INST_A2F_R_5_0 (.IN_IBUF(tcdm_rdata_p0[12]),.OUT_IBUF(tcdm_rdata_p0_int[12]));

	qlIBUF QL_INST_A2F_R_5_1 (.IN_IBUF(tcdm_rdata_p0[13]),.OUT_IBUF(tcdm_rdata_p0_int[13]));

	qlIBUF QL_INST_A2F_R_5_2 (.IN_IBUF(tcdm_rdata_p0[14]),.OUT_IBUF(tcdm_rdata_p0_int[14]));

	qlIBUF QL_INST_A2F_R_5_3 (.IN_IBUF(tcdm_rdata_p0[15]),.OUT_IBUF(tcdm_rdata_p0_int[15]));

	qlOBUF QL_INST_F2A_R_6_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[16]),.OUT_OBUF(tcdm_wdata_p0[16]));

	qlOBUF QL_INST_F2A_R_6_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[17]),.OUT_OBUF(tcdm_wdata_p0[17]));

	qlOBUF QL_INST_F2A_R_6_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[18]),.OUT_OBUF(tcdm_wdata_p0[18]));

	qlOBUF QL_INST_F2A_R_6_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[19]),.OUT_OBUF(tcdm_wdata_p0[19]));

	qlOBUF QL_INST_F2A_R_6_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[20]),.OUT_OBUF(tcdm_wdata_p0[20]));

	qlOBUF QL_INST_F2A_R_6_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[21]),.OUT_OBUF(tcdm_wdata_p0[21]));

	qlOBUF QL_INST_F2A_R_6_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[22]),.OUT_OBUF(tcdm_wdata_p0[22]));

	qlOBUF QL_INST_F2A_R_6_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[23]),.OUT_OBUF(tcdm_wdata_p0[23]));

	qlOBUF QL_INST_F2A_R_6_12 (.IN_OBUF(tcdm_addr_p0_dup_0[14]),.OUT_OBUF(tcdm_addr_p0[14]));

	qlOBUF QL_INST_F2A_R_6_13 (.IN_OBUF(tcdm_addr_p0_dup_0[15]),.OUT_OBUF(tcdm_addr_p0[15]));

	qlOBUF QL_INST_F2A_R_6_14 (.IN_OBUF(tcdm_addr_p0_dup_0[16]),.OUT_OBUF(tcdm_addr_p0[16]));

	qlOBUF QL_INST_F2A_R_6_15 (.IN_OBUF(tcdm_addr_p0_dup_0[17]),.OUT_OBUF(tcdm_addr_p0[17]));

	qlOBUF QL_INST_F2A_R_6_16 (.IN_OBUF(tcdm_addr_p0_dup_0[18]),.OUT_OBUF(tcdm_addr_p0[18]));

	qlOBUF QL_INST_F2A_R_6_17 (.IN_OBUF(tcdm_addr_p0_dup_0[19]),.OUT_OBUF(tcdm_addr_p0[19]));

	qlIBUF QL_INST_A2F_R_6_0 (.IN_IBUF(RESET[0]),.OUT_IBUF(RESET_int[0]));

	qlIBUF QL_INST_A2F_R_6_1 (.IN_IBUF(tcdm_rdata_p0[16]),.OUT_IBUF(tcdm_rdata_p0_int[16]));

	qlIBUF QL_INST_A2F_R_6_2 (.IN_IBUF(tcdm_rdata_p0[17]),.OUT_IBUF(tcdm_rdata_p0_int[17]));

	qlIBUF QL_INST_A2F_R_6_3 (.IN_IBUF(tcdm_rdata_p0[18]),.OUT_IBUF(tcdm_rdata_p0_int[18]));

	qlIBUF QL_INST_A2F_R_6_4 (.IN_IBUF(tcdm_rdata_p0[19]),.OUT_IBUF(tcdm_rdata_p0_int[19]));

	qlIBUF QL_INST_A2F_R_6_5 (.IN_IBUF(tcdm_rdata_p0[20]),.OUT_IBUF(tcdm_rdata_p0_int[20]));

	qlIBUF QL_INST_A2F_R_6_6 (.IN_IBUF(tcdm_rdata_p0[21]),.OUT_IBUF(tcdm_rdata_p0_int[21]));

	qlOBUF QL_INST_F2A_R_7_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[24]),.OUT_OBUF(tcdm_wdata_p0[24]));

	qlOBUF QL_INST_F2A_R_7_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[25]),.OUT_OBUF(tcdm_wdata_p0[25]));

	qlOBUF QL_INST_F2A_R_7_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[26]),.OUT_OBUF(tcdm_wdata_p0[26]));

	qlOBUF QL_INST_F2A_R_7_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[27]),.OUT_OBUF(tcdm_wdata_p0[27]));

	qlOBUF QL_INST_F2A_R_7_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[28]),.OUT_OBUF(tcdm_wdata_p0[28]));

	qlOBUF QL_INST_F2A_R_7_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[29]),.OUT_OBUF(tcdm_wdata_p0[29]));

	qlOBUF QL_INST_F2A_R_7_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[30]),.OUT_OBUF(tcdm_wdata_p0[30]));

	qlOBUF QL_INST_F2A_R_7_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[31]),.OUT_OBUF(tcdm_wdata_p0[31]));

	qlIBUF QL_INST_A2F_R_7_0 (.IN_IBUF(tcdm_rdata_p0[22]),.OUT_IBUF(tcdm_rdata_p0_int[22]));

	qlIBUF QL_INST_A2F_R_7_1 (.IN_IBUF(tcdm_rdata_p0[23]),.OUT_IBUF(tcdm_rdata_p0_int[23]));

	qlIBUF QL_INST_A2F_R_7_2 (.IN_IBUF(tcdm_rdata_p0[24]),.OUT_IBUF(tcdm_rdata_p0_int[24]));

	qlIBUF QL_INST_A2F_R_7_3 (.IN_IBUF(tcdm_rdata_p0[25]),.OUT_IBUF(tcdm_rdata_p0_int[25]));

	qlIBUF QL_INST_A2F_R_7_4 (.IN_IBUF(tcdm_rdata_p0[26]),.OUT_IBUF(tcdm_rdata_p0_int[26]));

	qlIBUF QL_INST_A2F_R_7_5 (.IN_IBUF(tcdm_rdata_p0[27]),.OUT_IBUF(tcdm_rdata_p0_int[27]));

	qlIBUF QL_INST_A2F_R_8_0 (.IN_IBUF(tcdm_rdata_p0[28]),.OUT_IBUF(tcdm_rdata_p0_int[28]));

	qlIBUF QL_INST_A2F_R_8_1 (.IN_IBUF(tcdm_rdata_p0[29]),.OUT_IBUF(tcdm_rdata_p0_int[29]));

	qlIBUF QL_INST_A2F_R_8_2 (.IN_IBUF(tcdm_rdata_p0[30]),.OUT_IBUF(tcdm_rdata_p0_int[30]));

	qlIBUF QL_INST_A2F_R_8_3 (.IN_IBUF(tcdm_rdata_p0[31]),.OUT_IBUF(tcdm_rdata_p0_int[31]));

	qlOBUF QL_INST_F2A_R_9_0 (.IN_OBUF(CLK_int_0__CAND0_TRSBR_33_padClk),.OUT_OBUF(tcdm_clk_p1));

	qlOBUF QL_INST_F2A_R_9_1 (.IN_OBUF(tcdm_req_p1_dup_0),.OUT_OBUF(tcdm_req_p1));

	qlOBUF QL_INST_F2A_R_9_2 (.IN_OBUF(tcdm_we_p1_dup_0),.OUT_OBUF(tcdm_we_p1));

	qlOBUF QL_INST_F2A_R_9_3 (.IN_OBUF(tcdm_be_p1_dup_0[0]),.OUT_OBUF(tcdm_be_p1[0]));

	qlOBUF QL_INST_F2A_R_9_4 (.IN_OBUF(tcdm_be_p1_dup_0[1]),.OUT_OBUF(tcdm_be_p1[1]));

	qlOBUF QL_INST_F2A_R_9_5 (.IN_OBUF(tcdm_be_p1_dup_0[2]),.OUT_OBUF(tcdm_be_p1[2]));

	qlOBUF QL_INST_F2A_R_9_6 (.IN_OBUF(tcdm_be_p1_dup_0[3]),.OUT_OBUF(tcdm_be_p1[3]));

	qlOBUF QL_INST_F2A_R_9_8 (.IN_OBUF(tcdm_addr_p1_dup_0[0]),.OUT_OBUF(tcdm_addr_p1[0]));

	qlOBUF QL_INST_F2A_R_9_9 (.IN_OBUF(tcdm_addr_p1_dup_0[1]),.OUT_OBUF(tcdm_addr_p1[1]));

	qlOBUF QL_INST_F2A_R_9_10 (.IN_OBUF(tcdm_addr_p1_dup_0[2]),.OUT_OBUF(tcdm_addr_p1[2]));

	qlOBUF QL_INST_F2A_R_9_11 (.IN_OBUF(tcdm_addr_p1_dup_0[3]),.OUT_OBUF(tcdm_addr_p1[3]));

	qlIBUF QL_INST_A2F_R_9_0 (.IN_IBUF(tcdm_rdata_p1[0]),.OUT_IBUF(tcdm_rdata_p1_int[0]));

	qlIBUF QL_INST_A2F_R_9_1 (.IN_IBUF(tcdm_rdata_p1[1]),.OUT_IBUF(tcdm_rdata_p1_int[1]));

	qlIBUF QL_INST_A2F_R_9_2 (.IN_IBUF(tcdm_rdata_p1[2]),.OUT_IBUF(tcdm_rdata_p1_int[2]));

	qlIBUF QL_INST_A2F_R_9_3 (.IN_IBUF(tcdm_rdata_p1[3]),.OUT_IBUF(tcdm_rdata_p1_int[3]));

	qlIBUF QL_INST_A2F_R_9_4 (.IN_IBUF(tcdm_valid_p1),.OUT_IBUF(tcdm_valid_p1_int));

	qlIBUF QL_INST_A2F_R_9_5 (.IN_IBUF(tcdm_gnt_p1),.OUT_IBUF(tcdm_gnt_p1_int));

	qlOBUF QL_INST_F2A_R_10_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[0]),.OUT_OBUF(tcdm_wdata_p1[0]));

	qlOBUF QL_INST_F2A_R_10_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[1]),.OUT_OBUF(tcdm_wdata_p1[1]));

	qlOBUF QL_INST_F2A_R_10_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[2]),.OUT_OBUF(tcdm_wdata_p1[2]));

	qlOBUF QL_INST_F2A_R_10_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[3]),.OUT_OBUF(tcdm_wdata_p1[3]));

	qlOBUF QL_INST_F2A_R_10_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[4]),.OUT_OBUF(tcdm_wdata_p1[4]));

	qlOBUF QL_INST_F2A_R_10_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[5]),.OUT_OBUF(tcdm_wdata_p1[5]));

	qlOBUF QL_INST_F2A_R_10_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[6]),.OUT_OBUF(tcdm_wdata_p1[6]));

	qlOBUF QL_INST_F2A_R_10_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[7]),.OUT_OBUF(tcdm_wdata_p1[7]));

	qlOBUF QL_INST_F2A_R_10_9 (.IN_OBUF(tcdm_addr_p1_dup_0[4]),.OUT_OBUF(tcdm_addr_p1[4]));

	qlOBUF QL_INST_F2A_R_10_10 (.IN_OBUF(tcdm_addr_p1_dup_0[5]),.OUT_OBUF(tcdm_addr_p1[5]));

	qlOBUF QL_INST_F2A_R_10_11 (.IN_OBUF(tcdm_addr_p1_dup_0[6]),.OUT_OBUF(tcdm_addr_p1[6]));

	qlOBUF QL_INST_F2A_R_10_12 (.IN_OBUF(tcdm_addr_p1_dup_0[7]),.OUT_OBUF(tcdm_addr_p1[7]));

	qlOBUF QL_INST_F2A_R_10_13 (.IN_OBUF(tcdm_addr_p1_dup_0[8]),.OUT_OBUF(tcdm_addr_p1[8]));

	qlOBUF QL_INST_F2A_R_10_14 (.IN_OBUF(tcdm_addr_p1_dup_0[9]),.OUT_OBUF(tcdm_addr_p1[9]));

	qlIBUF QL_INST_A2F_R_10_0 (.IN_IBUF(tcdm_rdata_p1[4]),.OUT_IBUF(tcdm_rdata_p1_int[4]));

	qlIBUF QL_INST_A2F_R_10_1 (.IN_IBUF(tcdm_rdata_p1[5]),.OUT_IBUF(tcdm_rdata_p1_int[5]));

	qlIBUF QL_INST_A2F_R_10_2 (.IN_IBUF(tcdm_rdata_p1[6]),.OUT_IBUF(tcdm_rdata_p1_int[6]));

	qlIBUF QL_INST_A2F_R_10_3 (.IN_IBUF(tcdm_rdata_p1[7]),.OUT_IBUF(tcdm_rdata_p1_int[7]));

	qlIBUF QL_INST_A2F_R_10_4 (.IN_IBUF(tcdm_rdata_p1[8]),.OUT_IBUF(tcdm_rdata_p1_int[8]));

	qlIBUF QL_INST_A2F_R_10_5 (.IN_IBUF(tcdm_rdata_p1[9]),.OUT_IBUF(tcdm_rdata_p1_int[9]));

	qlIBUF QL_INST_A2F_R_10_6 (.IN_IBUF(tcdm_rdata_p1[10]),.OUT_IBUF(tcdm_rdata_p1_int[10]));

	qlIBUF QL_INST_A2F_R_10_7 (.IN_IBUF(tcdm_rdata_p1[11]),.OUT_IBUF(tcdm_rdata_p1_int[11]));

	qlOBUF QL_INST_F2A_R_11_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[8]),.OUT_OBUF(tcdm_wdata_p1[8]));

	qlOBUF QL_INST_F2A_R_11_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[9]),.OUT_OBUF(tcdm_wdata_p1[9]));

	qlOBUF QL_INST_F2A_R_11_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[10]),.OUT_OBUF(tcdm_wdata_p1[10]));

	qlOBUF QL_INST_F2A_R_11_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[11]),.OUT_OBUF(tcdm_wdata_p1[11]));

	qlOBUF QL_INST_F2A_R_11_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[12]),.OUT_OBUF(tcdm_wdata_p1[12]));

	qlOBUF QL_INST_F2A_R_11_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[13]),.OUT_OBUF(tcdm_wdata_p1[13]));

	qlOBUF QL_INST_F2A_R_11_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[14]),.OUT_OBUF(tcdm_wdata_p1[14]));

	qlOBUF QL_INST_F2A_R_11_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[15]),.OUT_OBUF(tcdm_wdata_p1[15]));

	qlOBUF QL_INST_F2A_R_11_8 (.IN_OBUF(tcdm_addr_p1_dup_0[10]),.OUT_OBUF(tcdm_addr_p1[10]));

	qlOBUF QL_INST_F2A_R_11_9 (.IN_OBUF(tcdm_addr_p1_dup_0[11]),.OUT_OBUF(tcdm_addr_p1[11]));

	qlOBUF QL_INST_F2A_R_11_10 (.IN_OBUF(tcdm_addr_p1_dup_0[12]),.OUT_OBUF(tcdm_addr_p1[12]));

	qlOBUF QL_INST_F2A_R_11_11 (.IN_OBUF(tcdm_addr_p1_dup_0[13]),.OUT_OBUF(tcdm_addr_p1[13]));

	qlIBUF QL_INST_A2F_R_11_0 (.IN_IBUF(tcdm_rdata_p1[12]),.OUT_IBUF(tcdm_rdata_p1_int[12]));

	qlIBUF QL_INST_A2F_R_11_1 (.IN_IBUF(tcdm_rdata_p1[13]),.OUT_IBUF(tcdm_rdata_p1_int[13]));

	qlIBUF QL_INST_A2F_R_11_2 (.IN_IBUF(tcdm_rdata_p1[14]),.OUT_IBUF(tcdm_rdata_p1_int[14]));

	qlIBUF QL_INST_A2F_R_11_3 (.IN_IBUF(tcdm_rdata_p1[15]),.OUT_IBUF(tcdm_rdata_p1_int[15]));

	qlOBUF QL_INST_F2A_R_12_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[16]),.OUT_OBUF(tcdm_wdata_p1[16]));

	qlOBUF QL_INST_F2A_R_12_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[17]),.OUT_OBUF(tcdm_wdata_p1[17]));

	qlOBUF QL_INST_F2A_R_12_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[18]),.OUT_OBUF(tcdm_wdata_p1[18]));

	qlOBUF QL_INST_F2A_R_12_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[19]),.OUT_OBUF(tcdm_wdata_p1[19]));

	qlOBUF QL_INST_F2A_R_12_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[20]),.OUT_OBUF(tcdm_wdata_p1[20]));

	qlOBUF QL_INST_F2A_R_12_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[21]),.OUT_OBUF(tcdm_wdata_p1[21]));

	qlOBUF QL_INST_F2A_R_12_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[22]),.OUT_OBUF(tcdm_wdata_p1[22]));

	qlOBUF QL_INST_F2A_R_12_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[23]),.OUT_OBUF(tcdm_wdata_p1[23]));

	qlOBUF QL_INST_F2A_R_12_12 (.IN_OBUF(tcdm_addr_p1_dup_0[14]),.OUT_OBUF(tcdm_addr_p1[14]));

	qlOBUF QL_INST_F2A_R_12_13 (.IN_OBUF(tcdm_addr_p1_dup_0[15]),.OUT_OBUF(tcdm_addr_p1[15]));

	qlOBUF QL_INST_F2A_R_12_14 (.IN_OBUF(tcdm_addr_p1_dup_0[16]),.OUT_OBUF(tcdm_addr_p1[16]));

	qlOBUF QL_INST_F2A_R_12_15 (.IN_OBUF(tcdm_addr_p1_dup_0[17]),.OUT_OBUF(tcdm_addr_p1[17]));

	qlOBUF QL_INST_F2A_R_12_16 (.IN_OBUF(tcdm_addr_p1_dup_0[18]),.OUT_OBUF(tcdm_addr_p1[18]));

	qlOBUF QL_INST_F2A_R_12_17 (.IN_OBUF(tcdm_addr_p1_dup_0[19]),.OUT_OBUF(tcdm_addr_p1[19]));

	qlIBUF QL_INST_A2F_R_12_1 (.IN_IBUF(tcdm_rdata_p1[16]),.OUT_IBUF(tcdm_rdata_p1_int[16]));

	qlIBUF QL_INST_A2F_R_12_2 (.IN_IBUF(tcdm_rdata_p1[17]),.OUT_IBUF(tcdm_rdata_p1_int[17]));

	qlIBUF QL_INST_A2F_R_12_3 (.IN_IBUF(tcdm_rdata_p1[18]),.OUT_IBUF(tcdm_rdata_p1_int[18]));

	qlIBUF QL_INST_A2F_R_12_4 (.IN_IBUF(tcdm_rdata_p1[19]),.OUT_IBUF(tcdm_rdata_p1_int[19]));

	qlIBUF QL_INST_A2F_R_12_5 (.IN_IBUF(tcdm_rdata_p1[20]),.OUT_IBUF(tcdm_rdata_p1_int[20]));

	qlIBUF QL_INST_A2F_R_12_6 (.IN_IBUF(tcdm_rdata_p1[21]),.OUT_IBUF(tcdm_rdata_p1_int[21]));

	qlOBUF QL_INST_F2A_R_13_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[24]),.OUT_OBUF(tcdm_wdata_p1[24]));

	qlOBUF QL_INST_F2A_R_13_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[25]),.OUT_OBUF(tcdm_wdata_p1[25]));

	qlOBUF QL_INST_F2A_R_13_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[26]),.OUT_OBUF(tcdm_wdata_p1[26]));

	qlOBUF QL_INST_F2A_R_13_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[27]),.OUT_OBUF(tcdm_wdata_p1[27]));

	qlOBUF QL_INST_F2A_R_13_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[28]),.OUT_OBUF(tcdm_wdata_p1[28]));

	qlOBUF QL_INST_F2A_R_13_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[29]),.OUT_OBUF(tcdm_wdata_p1[29]));

	qlOBUF QL_INST_F2A_R_13_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[30]),.OUT_OBUF(tcdm_wdata_p1[30]));

	qlOBUF QL_INST_F2A_R_13_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[31]),.OUT_OBUF(tcdm_wdata_p1[31]));

	qlIBUF QL_INST_A2F_R_13_0 (.IN_IBUF(tcdm_rdata_p1[22]),.OUT_IBUF(tcdm_rdata_p1_int[22]));

	qlIBUF QL_INST_A2F_R_13_1 (.IN_IBUF(tcdm_rdata_p1[23]),.OUT_IBUF(tcdm_rdata_p1_int[23]));

	qlIBUF QL_INST_A2F_R_13_2 (.IN_IBUF(tcdm_rdata_p1[24]),.OUT_IBUF(tcdm_rdata_p1_int[24]));

	qlIBUF QL_INST_A2F_R_13_3 (.IN_IBUF(tcdm_rdata_p1[25]),.OUT_IBUF(tcdm_rdata_p1_int[25]));

	qlIBUF QL_INST_A2F_R_13_4 (.IN_IBUF(tcdm_rdata_p1[26]),.OUT_IBUF(tcdm_rdata_p1_int[26]));

	qlIBUF QL_INST_A2F_R_13_5 (.IN_IBUF(tcdm_rdata_p1[27]),.OUT_IBUF(tcdm_rdata_p1_int[27]));

	qlIBUF QL_INST_A2F_R_14_0 (.IN_IBUF(tcdm_rdata_p1[28]),.OUT_IBUF(tcdm_rdata_p1_int[28]));

	qlIBUF QL_INST_A2F_R_14_1 (.IN_IBUF(tcdm_rdata_p1[29]),.OUT_IBUF(tcdm_rdata_p1_int[29]));

	qlIBUF QL_INST_A2F_R_14_2 (.IN_IBUF(tcdm_rdata_p1[30]),.OUT_IBUF(tcdm_rdata_p1_int[30]));

	qlIBUF QL_INST_A2F_R_14_3 (.IN_IBUF(tcdm_rdata_p1[31]),.OUT_IBUF(tcdm_rdata_p1_int[31]));

	qlOBUF QL_INST_F2A_R_17_0 (.IN_OBUF(CLK_int_0__CAND0_BRSTR_33_padClk),.OUT_OBUF(tcdm_clk_p2));

	qlOBUF QL_INST_F2A_R_17_1 (.IN_OBUF(tcdm_req_p2_dup_0),.OUT_OBUF(tcdm_req_p2));

	qlOBUF QL_INST_F2A_R_17_2 (.IN_OBUF(tcdm_we_p2_dup_0),.OUT_OBUF(tcdm_we_p2));

	qlOBUF QL_INST_F2A_R_17_3 (.IN_OBUF(tcdm_be_p2_dup_0[0]),.OUT_OBUF(tcdm_be_p2[0]));

	qlOBUF QL_INST_F2A_R_17_4 (.IN_OBUF(tcdm_be_p2_dup_0[1]),.OUT_OBUF(tcdm_be_p2[1]));

	qlOBUF QL_INST_F2A_R_17_5 (.IN_OBUF(tcdm_be_p2_dup_0[2]),.OUT_OBUF(tcdm_be_p2[2]));

	qlOBUF QL_INST_F2A_R_17_6 (.IN_OBUF(tcdm_be_p2_dup_0[3]),.OUT_OBUF(tcdm_be_p2[3]));

	qlOBUF QL_INST_F2A_R_17_8 (.IN_OBUF(tcdm_addr_p2_dup_0[0]),.OUT_OBUF(tcdm_addr_p2[0]));

	qlOBUF QL_INST_F2A_R_17_9 (.IN_OBUF(tcdm_addr_p2_dup_0[1]),.OUT_OBUF(tcdm_addr_p2[1]));

	qlOBUF QL_INST_F2A_R_17_10 (.IN_OBUF(tcdm_addr_p2_dup_0[2]),.OUT_OBUF(tcdm_addr_p2[2]));

	qlOBUF QL_INST_F2A_R_17_11 (.IN_OBUF(tcdm_addr_p2_dup_0[3]),.OUT_OBUF(tcdm_addr_p2[3]));

	qlIBUF QL_INST_A2F_R_17_0 (.IN_IBUF(tcdm_rdata_p2[0]),.OUT_IBUF(tcdm_rdata_p2_int[0]));

	qlIBUF QL_INST_A2F_R_17_1 (.IN_IBUF(tcdm_rdata_p2[1]),.OUT_IBUF(tcdm_rdata_p2_int[1]));

	qlIBUF QL_INST_A2F_R_17_2 (.IN_IBUF(tcdm_rdata_p2[2]),.OUT_IBUF(tcdm_rdata_p2_int[2]));

	qlIBUF QL_INST_A2F_R_17_3 (.IN_IBUF(tcdm_rdata_p2[3]),.OUT_IBUF(tcdm_rdata_p2_int[3]));

	qlIBUF QL_INST_A2F_R_17_4 (.IN_IBUF(tcdm_valid_p2),.OUT_IBUF(tcdm_valid_p2_int));

	qlIBUF QL_INST_A2F_R_17_5 (.IN_IBUF(tcdm_gnt_p2),.OUT_IBUF(tcdm_gnt_p2_int));

	qlOBUF QL_INST_F2A_R_18_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[0]),.OUT_OBUF(tcdm_wdata_p2[0]));

	qlOBUF QL_INST_F2A_R_18_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[1]),.OUT_OBUF(tcdm_wdata_p2[1]));

	qlOBUF QL_INST_F2A_R_18_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[2]),.OUT_OBUF(tcdm_wdata_p2[2]));

	qlOBUF QL_INST_F2A_R_18_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[3]),.OUT_OBUF(tcdm_wdata_p2[3]));

	qlOBUF QL_INST_F2A_R_18_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[4]),.OUT_OBUF(tcdm_wdata_p2[4]));

	qlOBUF QL_INST_F2A_R_18_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[5]),.OUT_OBUF(tcdm_wdata_p2[5]));

	qlOBUF QL_INST_F2A_R_18_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[6]),.OUT_OBUF(tcdm_wdata_p2[6]));

	qlOBUF QL_INST_F2A_R_18_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[7]),.OUT_OBUF(tcdm_wdata_p2[7]));

	qlOBUF QL_INST_F2A_R_18_9 (.IN_OBUF(tcdm_addr_p2_dup_0[4]),.OUT_OBUF(tcdm_addr_p2[4]));

	qlOBUF QL_INST_F2A_R_18_10 (.IN_OBUF(tcdm_addr_p2_dup_0[5]),.OUT_OBUF(tcdm_addr_p2[5]));

	qlOBUF QL_INST_F2A_R_18_11 (.IN_OBUF(tcdm_addr_p2_dup_0[6]),.OUT_OBUF(tcdm_addr_p2[6]));

	qlOBUF QL_INST_F2A_R_18_12 (.IN_OBUF(tcdm_addr_p2_dup_0[7]),.OUT_OBUF(tcdm_addr_p2[7]));

	qlOBUF QL_INST_F2A_R_18_13 (.IN_OBUF(tcdm_addr_p2_dup_0[8]),.OUT_OBUF(tcdm_addr_p2[8]));

	qlOBUF QL_INST_F2A_R_18_14 (.IN_OBUF(tcdm_addr_p2_dup_0[9]),.OUT_OBUF(tcdm_addr_p2[9]));

	qlIBUF QL_INST_A2F_R_18_0 (.IN_IBUF(tcdm_rdata_p2[4]),.OUT_IBUF(tcdm_rdata_p2_int[4]));

	qlIBUF QL_INST_A2F_R_18_1 (.IN_IBUF(tcdm_rdata_p2[5]),.OUT_IBUF(tcdm_rdata_p2_int[5]));

	qlIBUF QL_INST_A2F_R_18_2 (.IN_IBUF(tcdm_rdata_p2[6]),.OUT_IBUF(tcdm_rdata_p2_int[6]));

	qlIBUF QL_INST_A2F_R_18_3 (.IN_IBUF(tcdm_rdata_p2[7]),.OUT_IBUF(tcdm_rdata_p2_int[7]));

	qlIBUF QL_INST_A2F_R_18_4 (.IN_IBUF(tcdm_rdata_p2[8]),.OUT_IBUF(tcdm_rdata_p2_int[8]));

	qlIBUF QL_INST_A2F_R_18_5 (.IN_IBUF(tcdm_rdata_p2[9]),.OUT_IBUF(tcdm_rdata_p2_int[9]));

	qlIBUF QL_INST_A2F_R_18_6 (.IN_IBUF(tcdm_rdata_p2[10]),.OUT_IBUF(tcdm_rdata_p2_int[10]));

	qlIBUF QL_INST_A2F_R_18_7 (.IN_IBUF(tcdm_rdata_p2[11]),.OUT_IBUF(tcdm_rdata_p2_int[11]));

	qlOBUF QL_INST_F2A_R_19_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[8]),.OUT_OBUF(tcdm_wdata_p2[8]));

	qlOBUF QL_INST_F2A_R_19_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[9]),.OUT_OBUF(tcdm_wdata_p2[9]));

	qlOBUF QL_INST_F2A_R_19_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[10]),.OUT_OBUF(tcdm_wdata_p2[10]));

	qlOBUF QL_INST_F2A_R_19_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[11]),.OUT_OBUF(tcdm_wdata_p2[11]));

	qlOBUF QL_INST_F2A_R_19_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[12]),.OUT_OBUF(tcdm_wdata_p2[12]));

	qlOBUF QL_INST_F2A_R_19_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[13]),.OUT_OBUF(tcdm_wdata_p2[13]));

	qlOBUF QL_INST_F2A_R_19_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[14]),.OUT_OBUF(tcdm_wdata_p2[14]));

	qlOBUF QL_INST_F2A_R_19_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[15]),.OUT_OBUF(tcdm_wdata_p2[15]));

	qlOBUF QL_INST_F2A_R_19_8 (.IN_OBUF(tcdm_addr_p2_dup_0[10]),.OUT_OBUF(tcdm_addr_p2[10]));

	qlOBUF QL_INST_F2A_R_19_9 (.IN_OBUF(tcdm_addr_p2_dup_0[11]),.OUT_OBUF(tcdm_addr_p2[11]));

	qlOBUF QL_INST_F2A_R_19_10 (.IN_OBUF(tcdm_addr_p2_dup_0[12]),.OUT_OBUF(tcdm_addr_p2[12]));

	qlOBUF QL_INST_F2A_R_19_11 (.IN_OBUF(tcdm_addr_p2_dup_0[13]),.OUT_OBUF(tcdm_addr_p2[13]));

	qlIBUF QL_INST_A2F_R_19_0 (.IN_IBUF(tcdm_rdata_p2[12]),.OUT_IBUF(tcdm_rdata_p2_int[12]));

	qlIBUF QL_INST_A2F_R_19_1 (.IN_IBUF(tcdm_rdata_p2[13]),.OUT_IBUF(tcdm_rdata_p2_int[13]));

	qlIBUF QL_INST_A2F_R_19_2 (.IN_IBUF(tcdm_rdata_p2[14]),.OUT_IBUF(tcdm_rdata_p2_int[14]));

	qlIBUF QL_INST_A2F_R_19_3 (.IN_IBUF(tcdm_rdata_p2[15]),.OUT_IBUF(tcdm_rdata_p2_int[15]));

	qlOBUF QL_INST_F2A_R_20_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[16]),.OUT_OBUF(tcdm_wdata_p2[16]));

	qlOBUF QL_INST_F2A_R_20_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[17]),.OUT_OBUF(tcdm_wdata_p2[17]));

	qlOBUF QL_INST_F2A_R_20_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[18]),.OUT_OBUF(tcdm_wdata_p2[18]));

	qlOBUF QL_INST_F2A_R_20_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[19]),.OUT_OBUF(tcdm_wdata_p2[19]));

	qlOBUF QL_INST_F2A_R_20_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[20]),.OUT_OBUF(tcdm_wdata_p2[20]));

	qlOBUF QL_INST_F2A_R_20_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[21]),.OUT_OBUF(tcdm_wdata_p2[21]));

	qlOBUF QL_INST_F2A_R_20_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[22]),.OUT_OBUF(tcdm_wdata_p2[22]));

	qlOBUF QL_INST_F2A_R_20_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[23]),.OUT_OBUF(tcdm_wdata_p2[23]));

	qlOBUF QL_INST_F2A_R_20_12 (.IN_OBUF(tcdm_addr_p2_dup_0[14]),.OUT_OBUF(tcdm_addr_p2[14]));

	qlOBUF QL_INST_F2A_R_20_13 (.IN_OBUF(tcdm_addr_p2_dup_0[15]),.OUT_OBUF(tcdm_addr_p2[15]));

	qlOBUF QL_INST_F2A_R_20_14 (.IN_OBUF(tcdm_addr_p2_dup_0[16]),.OUT_OBUF(tcdm_addr_p2[16]));

	qlOBUF QL_INST_F2A_R_20_15 (.IN_OBUF(tcdm_addr_p2_dup_0[17]),.OUT_OBUF(tcdm_addr_p2[17]));

	qlOBUF QL_INST_F2A_R_20_16 (.IN_OBUF(tcdm_addr_p2_dup_0[18]),.OUT_OBUF(tcdm_addr_p2[18]));

	qlOBUF QL_INST_F2A_R_20_17 (.IN_OBUF(tcdm_addr_p2_dup_0[19]),.OUT_OBUF(tcdm_addr_p2[19]));

	qlIBUF QL_INST_A2F_R_20_1 (.IN_IBUF(tcdm_rdata_p2[16]),.OUT_IBUF(tcdm_rdata_p2_int[16]));

	qlIBUF QL_INST_A2F_R_20_2 (.IN_IBUF(tcdm_rdata_p2[17]),.OUT_IBUF(tcdm_rdata_p2_int[17]));

	qlIBUF QL_INST_A2F_R_20_3 (.IN_IBUF(tcdm_rdata_p2[18]),.OUT_IBUF(tcdm_rdata_p2_int[18]));

	qlIBUF QL_INST_A2F_R_20_4 (.IN_IBUF(tcdm_rdata_p2[19]),.OUT_IBUF(tcdm_rdata_p2_int[19]));

	qlIBUF QL_INST_A2F_R_20_5 (.IN_IBUF(tcdm_rdata_p2[20]),.OUT_IBUF(tcdm_rdata_p2_int[20]));

	qlIBUF QL_INST_A2F_R_20_6 (.IN_IBUF(tcdm_rdata_p2[21]),.OUT_IBUF(tcdm_rdata_p2_int[21]));

	qlOBUF QL_INST_F2A_R_21_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[24]),.OUT_OBUF(tcdm_wdata_p2[24]));

	qlOBUF QL_INST_F2A_R_21_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[25]),.OUT_OBUF(tcdm_wdata_p2[25]));

	qlOBUF QL_INST_F2A_R_21_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[26]),.OUT_OBUF(tcdm_wdata_p2[26]));

	qlOBUF QL_INST_F2A_R_21_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[27]),.OUT_OBUF(tcdm_wdata_p2[27]));

	qlOBUF QL_INST_F2A_R_21_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[28]),.OUT_OBUF(tcdm_wdata_p2[28]));

	qlOBUF QL_INST_F2A_R_21_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[29]),.OUT_OBUF(tcdm_wdata_p2[29]));

	qlOBUF QL_INST_F2A_R_21_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[30]),.OUT_OBUF(tcdm_wdata_p2[30]));

	qlOBUF QL_INST_F2A_R_21_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[31]),.OUT_OBUF(tcdm_wdata_p2[31]));

	qlIBUF QL_INST_A2F_R_21_0 (.IN_IBUF(tcdm_rdata_p2[22]),.OUT_IBUF(tcdm_rdata_p2_int[22]));

	qlIBUF QL_INST_A2F_R_21_1 (.IN_IBUF(tcdm_rdata_p2[23]),.OUT_IBUF(tcdm_rdata_p2_int[23]));

	qlIBUF QL_INST_A2F_R_21_2 (.IN_IBUF(tcdm_rdata_p2[24]),.OUT_IBUF(tcdm_rdata_p2_int[24]));

	qlIBUF QL_INST_A2F_R_21_3 (.IN_IBUF(tcdm_rdata_p2[25]),.OUT_IBUF(tcdm_rdata_p2_int[25]));

	qlIBUF QL_INST_A2F_R_21_4 (.IN_IBUF(tcdm_rdata_p2[26]),.OUT_IBUF(tcdm_rdata_p2_int[26]));

	qlIBUF QL_INST_A2F_R_21_5 (.IN_IBUF(tcdm_rdata_p2[27]),.OUT_IBUF(tcdm_rdata_p2_int[27]));

	qlIBUF QL_INST_A2F_R_22_0 (.IN_IBUF(tcdm_rdata_p2[28]),.OUT_IBUF(tcdm_rdata_p2_int[28]));

	qlIBUF QL_INST_A2F_R_22_1 (.IN_IBUF(tcdm_rdata_p2[29]),.OUT_IBUF(tcdm_rdata_p2_int[29]));

	qlIBUF QL_INST_A2F_R_22_2 (.IN_IBUF(tcdm_rdata_p2[30]),.OUT_IBUF(tcdm_rdata_p2_int[30]));

	qlIBUF QL_INST_A2F_R_22_3 (.IN_IBUF(tcdm_rdata_p2[31]),.OUT_IBUF(tcdm_rdata_p2_int[31]));

	qlOBUF QL_INST_F2A_R_23_0 (.IN_OBUF(CLK_int_0__CAND0_BRSTR_33_padClk),.OUT_OBUF(tcdm_clk_p3));

	qlOBUF QL_INST_F2A_R_23_1 (.IN_OBUF(tcdm_req_p3_dup_0),.OUT_OBUF(tcdm_req_p3));

	qlOBUF QL_INST_F2A_R_23_2 (.IN_OBUF(tcdm_we_p3_dup_0),.OUT_OBUF(tcdm_we_p3));

	qlOBUF QL_INST_F2A_R_23_3 (.IN_OBUF(tcdm_be_p3_dup_0[0]),.OUT_OBUF(tcdm_be_p3[0]));

	qlOBUF QL_INST_F2A_R_23_4 (.IN_OBUF(tcdm_be_p3_dup_0[1]),.OUT_OBUF(tcdm_be_p3[1]));

	qlOBUF QL_INST_F2A_R_23_5 (.IN_OBUF(tcdm_be_p3_dup_0[2]),.OUT_OBUF(tcdm_be_p3[2]));

	qlOBUF QL_INST_F2A_R_23_6 (.IN_OBUF(tcdm_be_p3_dup_0[3]),.OUT_OBUF(tcdm_be_p3[3]));

	qlOBUF QL_INST_F2A_R_23_8 (.IN_OBUF(tcdm_addr_p3_dup_0[0]),.OUT_OBUF(tcdm_addr_p3[0]));

	qlOBUF QL_INST_F2A_R_23_9 (.IN_OBUF(tcdm_addr_p3_dup_0[1]),.OUT_OBUF(tcdm_addr_p3[1]));

	qlOBUF QL_INST_F2A_R_23_10 (.IN_OBUF(tcdm_addr_p3_dup_0[2]),.OUT_OBUF(tcdm_addr_p3[2]));

	qlOBUF QL_INST_F2A_R_23_11 (.IN_OBUF(tcdm_addr_p3_dup_0[3]),.OUT_OBUF(tcdm_addr_p3[3]));

	qlIBUF QL_INST_A2F_R_23_0 (.IN_IBUF(tcdm_rdata_p3[0]),.OUT_IBUF(tcdm_rdata_p3_int[0]));

	qlIBUF QL_INST_A2F_R_23_1 (.IN_IBUF(tcdm_rdata_p3[1]),.OUT_IBUF(tcdm_rdata_p3_int[1]));

	qlIBUF QL_INST_A2F_R_23_2 (.IN_IBUF(tcdm_rdata_p3[2]),.OUT_IBUF(tcdm_rdata_p3_int[2]));

	qlIBUF QL_INST_A2F_R_23_3 (.IN_IBUF(tcdm_rdata_p3[3]),.OUT_IBUF(tcdm_rdata_p3_int[3]));

	qlIBUF QL_INST_A2F_R_23_4 (.IN_IBUF(tcdm_valid_p3),.OUT_IBUF(tcdm_valid_p3_int));

	qlIBUF QL_INST_A2F_R_23_5 (.IN_IBUF(tcdm_gnt_p3),.OUT_IBUF(tcdm_gnt_p3_int));

	qlOBUF QL_INST_F2A_R_24_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[0]),.OUT_OBUF(tcdm_wdata_p3[0]));

	qlOBUF QL_INST_F2A_R_24_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[1]),.OUT_OBUF(tcdm_wdata_p3[1]));

	qlOBUF QL_INST_F2A_R_24_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[2]),.OUT_OBUF(tcdm_wdata_p3[2]));

	qlOBUF QL_INST_F2A_R_24_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[3]),.OUT_OBUF(tcdm_wdata_p3[3]));

	qlOBUF QL_INST_F2A_R_24_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[5]),.OUT_OBUF(tcdm_wdata_p3[5]));

	qlOBUF QL_INST_F2A_R_24_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[4]),.OUT_OBUF(tcdm_wdata_p3[4]));

	qlOBUF QL_INST_F2A_R_24_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[6]),.OUT_OBUF(tcdm_wdata_p3[6]));

	qlOBUF QL_INST_F2A_R_24_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[7]),.OUT_OBUF(tcdm_wdata_p3[7]));

	qlOBUF QL_INST_F2A_R_24_9 (.IN_OBUF(tcdm_addr_p3_dup_0[4]),.OUT_OBUF(tcdm_addr_p3[4]));

	qlOBUF QL_INST_F2A_R_24_10 (.IN_OBUF(tcdm_addr_p3_dup_0[5]),.OUT_OBUF(tcdm_addr_p3[5]));

	qlOBUF QL_INST_F2A_R_24_11 (.IN_OBUF(tcdm_addr_p3_dup_0[6]),.OUT_OBUF(tcdm_addr_p3[6]));

	qlOBUF QL_INST_F2A_R_24_12 (.IN_OBUF(tcdm_addr_p3_dup_0[7]),.OUT_OBUF(tcdm_addr_p3[7]));

	qlOBUF QL_INST_F2A_R_24_13 (.IN_OBUF(tcdm_addr_p3_dup_0[8]),.OUT_OBUF(tcdm_addr_p3[8]));

	qlOBUF QL_INST_F2A_R_24_14 (.IN_OBUF(tcdm_addr_p3_dup_0[9]),.OUT_OBUF(tcdm_addr_p3[9]));

	qlIBUF QL_INST_A2F_R_24_0 (.IN_IBUF(tcdm_rdata_p3[4]),.OUT_IBUF(tcdm_rdata_p3_int[4]));

	qlIBUF QL_INST_A2F_R_24_1 (.IN_IBUF(tcdm_rdata_p3[5]),.OUT_IBUF(tcdm_rdata_p3_int[5]));

	qlIBUF QL_INST_A2F_R_24_2 (.IN_IBUF(tcdm_rdata_p3[6]),.OUT_IBUF(tcdm_rdata_p3_int[6]));

	qlIBUF QL_INST_A2F_R_24_3 (.IN_IBUF(tcdm_rdata_p3[7]),.OUT_IBUF(tcdm_rdata_p3_int[7]));

	qlIBUF QL_INST_A2F_R_24_4 (.IN_IBUF(tcdm_rdata_p3[8]),.OUT_IBUF(tcdm_rdata_p3_int[8]));

	qlIBUF QL_INST_A2F_R_24_5 (.IN_IBUF(tcdm_rdata_p3[9]),.OUT_IBUF(tcdm_rdata_p3_int[9]));

	qlIBUF QL_INST_A2F_R_24_6 (.IN_IBUF(tcdm_rdata_p3[10]),.OUT_IBUF(tcdm_rdata_p3_int[10]));

	qlIBUF QL_INST_A2F_R_24_7 (.IN_IBUF(tcdm_rdata_p3[11]),.OUT_IBUF(tcdm_rdata_p3_int[11]));

	qlOBUF QL_INST_F2A_R_25_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[8]),.OUT_OBUF(tcdm_wdata_p3[8]));

	qlOBUF QL_INST_F2A_R_25_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[9]),.OUT_OBUF(tcdm_wdata_p3[9]));

	qlOBUF QL_INST_F2A_R_25_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[10]),.OUT_OBUF(tcdm_wdata_p3[10]));

	qlOBUF QL_INST_F2A_R_25_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[11]),.OUT_OBUF(tcdm_wdata_p3[11]));

	qlOBUF QL_INST_F2A_R_25_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[12]),.OUT_OBUF(tcdm_wdata_p3[12]));

	qlOBUF QL_INST_F2A_R_25_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[13]),.OUT_OBUF(tcdm_wdata_p3[13]));

	qlOBUF QL_INST_F2A_R_25_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[14]),.OUT_OBUF(tcdm_wdata_p3[14]));

	qlOBUF QL_INST_F2A_R_25_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[15]),.OUT_OBUF(tcdm_wdata_p3[15]));

	qlOBUF QL_INST_F2A_R_25_8 (.IN_OBUF(tcdm_addr_p3_dup_0[10]),.OUT_OBUF(tcdm_addr_p3[10]));

	qlOBUF QL_INST_F2A_R_25_9 (.IN_OBUF(tcdm_addr_p3_dup_0[11]),.OUT_OBUF(tcdm_addr_p3[11]));

	qlOBUF QL_INST_F2A_R_25_10 (.IN_OBUF(tcdm_addr_p3_dup_0[12]),.OUT_OBUF(tcdm_addr_p3[12]));

	qlOBUF QL_INST_F2A_R_25_11 (.IN_OBUF(tcdm_addr_p3_dup_0[13]),.OUT_OBUF(tcdm_addr_p3[13]));

	qlIBUF QL_INST_A2F_R_25_0 (.IN_IBUF(tcdm_rdata_p3[12]),.OUT_IBUF(tcdm_rdata_p3_int[12]));

	qlIBUF QL_INST_A2F_R_25_1 (.IN_IBUF(tcdm_rdata_p3[13]),.OUT_IBUF(tcdm_rdata_p3_int[13]));

	qlIBUF QL_INST_A2F_R_25_2 (.IN_IBUF(tcdm_rdata_p3[14]),.OUT_IBUF(tcdm_rdata_p3_int[14]));

	qlIBUF QL_INST_A2F_R_25_3 (.IN_IBUF(tcdm_rdata_p3[15]),.OUT_IBUF(tcdm_rdata_p3_int[15]));

	qlOBUF QL_INST_F2A_R_26_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[16]),.OUT_OBUF(tcdm_wdata_p3[16]));

	qlOBUF QL_INST_F2A_R_26_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[17]),.OUT_OBUF(tcdm_wdata_p3[17]));

	qlOBUF QL_INST_F2A_R_26_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[18]),.OUT_OBUF(tcdm_wdata_p3[18]));

	qlOBUF QL_INST_F2A_R_26_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[19]),.OUT_OBUF(tcdm_wdata_p3[19]));

	qlOBUF QL_INST_F2A_R_26_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[20]),.OUT_OBUF(tcdm_wdata_p3[20]));

	qlOBUF QL_INST_F2A_R_26_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[21]),.OUT_OBUF(tcdm_wdata_p3[21]));

	qlOBUF QL_INST_F2A_R_26_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[22]),.OUT_OBUF(tcdm_wdata_p3[22]));

	qlOBUF QL_INST_F2A_R_26_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[23]),.OUT_OBUF(tcdm_wdata_p3[23]));

	qlOBUF QL_INST_F2A_R_26_12 (.IN_OBUF(tcdm_addr_p3_dup_0[14]),.OUT_OBUF(tcdm_addr_p3[14]));

	qlOBUF QL_INST_F2A_R_26_13 (.IN_OBUF(tcdm_addr_p3_dup_0[15]),.OUT_OBUF(tcdm_addr_p3[15]));

	qlOBUF QL_INST_F2A_R_26_14 (.IN_OBUF(tcdm_addr_p3_dup_0[16]),.OUT_OBUF(tcdm_addr_p3[16]));

	qlOBUF QL_INST_F2A_R_26_15 (.IN_OBUF(tcdm_addr_p3_dup_0[17]),.OUT_OBUF(tcdm_addr_p3[17]));

	qlOBUF QL_INST_F2A_R_26_16 (.IN_OBUF(tcdm_addr_p3_dup_0[18]),.OUT_OBUF(tcdm_addr_p3[18]));

	qlOBUF QL_INST_F2A_R_26_17 (.IN_OBUF(tcdm_addr_p3_dup_0[19]),.OUT_OBUF(tcdm_addr_p3[19]));

	qlIBUF QL_INST_A2F_R_26_1 (.IN_IBUF(tcdm_rdata_p3[16]),.OUT_IBUF(tcdm_rdata_p3_int[16]));

	qlIBUF QL_INST_A2F_R_26_2 (.IN_IBUF(tcdm_rdata_p3[17]),.OUT_IBUF(tcdm_rdata_p3_int[17]));

	qlIBUF QL_INST_A2F_R_26_3 (.IN_IBUF(tcdm_rdata_p3[18]),.OUT_IBUF(tcdm_rdata_p3_int[18]));

	qlIBUF QL_INST_A2F_R_26_4 (.IN_IBUF(tcdm_rdata_p3[19]),.OUT_IBUF(tcdm_rdata_p3_int[19]));

	qlIBUF QL_INST_A2F_R_26_5 (.IN_IBUF(tcdm_rdata_p3[20]),.OUT_IBUF(tcdm_rdata_p3_int[20]));

	qlIBUF QL_INST_A2F_R_26_6 (.IN_IBUF(tcdm_rdata_p3[21]),.OUT_IBUF(tcdm_rdata_p3_int[21]));

	qlOBUF QL_INST_F2A_R_27_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[24]),.OUT_OBUF(tcdm_wdata_p3[24]));

	qlOBUF QL_INST_F2A_R_27_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[25]),.OUT_OBUF(tcdm_wdata_p3[25]));

	qlOBUF QL_INST_F2A_R_27_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[26]),.OUT_OBUF(tcdm_wdata_p3[26]));

	qlOBUF QL_INST_F2A_R_27_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[27]),.OUT_OBUF(tcdm_wdata_p3[27]));

	qlOBUF QL_INST_F2A_R_27_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[28]),.OUT_OBUF(tcdm_wdata_p3[28]));

	qlOBUF QL_INST_F2A_R_27_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[29]),.OUT_OBUF(tcdm_wdata_p3[29]));

	qlOBUF QL_INST_F2A_R_27_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[30]),.OUT_OBUF(tcdm_wdata_p3[30]));

	qlOBUF QL_INST_F2A_R_27_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[31]),.OUT_OBUF(tcdm_wdata_p3[31]));

	qlIBUF QL_INST_A2F_R_27_0 (.IN_IBUF(tcdm_rdata_p3[22]),.OUT_IBUF(tcdm_rdata_p3_int[22]));

	qlIBUF QL_INST_A2F_R_27_1 (.IN_IBUF(tcdm_rdata_p3[23]),.OUT_IBUF(tcdm_rdata_p3_int[23]));

	qlIBUF QL_INST_A2F_R_27_2 (.IN_IBUF(tcdm_rdata_p3[24]),.OUT_IBUF(tcdm_rdata_p3_int[24]));

	qlIBUF QL_INST_A2F_R_27_3 (.IN_IBUF(tcdm_rdata_p3[25]),.OUT_IBUF(tcdm_rdata_p3_int[25]));

	qlIBUF QL_INST_A2F_R_27_4 (.IN_IBUF(tcdm_rdata_p3[26]),.OUT_IBUF(tcdm_rdata_p3_int[26]));

	qlIBUF QL_INST_A2F_R_27_5 (.IN_IBUF(tcdm_rdata_p3[27]),.OUT_IBUF(tcdm_rdata_p3_int[27]));

	qlIBUF QL_INST_A2F_R_28_0 (.IN_IBUF(tcdm_rdata_p3[28]),.OUT_IBUF(tcdm_rdata_p3_int[28]));

	qlIBUF QL_INST_A2F_R_28_1 (.IN_IBUF(tcdm_rdata_p3[29]),.OUT_IBUF(tcdm_rdata_p3_int[29]));

	qlIBUF QL_INST_A2F_R_28_2 (.IN_IBUF(tcdm_rdata_p3[30]),.OUT_IBUF(tcdm_rdata_p3_int[30]));

	qlIBUF QL_INST_A2F_R_28_3 (.IN_IBUF(tcdm_rdata_p3[31]),.OUT_IBUF(tcdm_rdata_p3_int[31]));

	qlIBUF QL_INST_A2F_R_29_2 (.IN_IBUF(RESET[1]),.OUT_IBUF(RESET_int[1]));

	qlIBUF QL_INST_A2F_B_3_2 (.IN_IBUF(m1_oper0_rdata[31]),.OUT_IBUF(m1_oper0_rdata_int[31]));

	qlIBUF QL_INST_A2F_B_3_3 (.IN_IBUF(m1_oper0_rdata[30]),.OUT_IBUF(m1_oper0_rdata_int[30]));

	qlIBUF QL_INST_A2F_B_3_4 (.IN_IBUF(m1_oper0_rdata[29]),.OUT_IBUF(m1_oper0_rdata_int[29]));

	qlIBUF QL_INST_A2F_B_3_5 (.IN_IBUF(m1_oper0_rdata[28]),.OUT_IBUF(m1_oper0_rdata_int[28]));

	qlOBUF QL_INST_F2A_B_4_0 (.IN_OBUF(CLK_int_0__CAND0_BLSBL_4_padClk),.OUT_OBUF(m1_oper0_wclk));

	qlOBUF QL_INST_F2A_B_4_2 (.IN_OBUF(m0_oper0_wmode_dup_0[1]),.OUT_OBUF(m1_oper0_wmode[1]));

	qlOBUF QL_INST_F2A_B_4_3 (.IN_OBUF(m0_oper0_wmode_dup_0[0]),.OUT_OBUF(m1_oper0_wmode[0]));

	qlOBUF QL_INST_F2A_B_4_4 (.IN_OBUF(m1_oper0_wdata_dup_0[31]),.OUT_OBUF(m1_oper0_wdata[31]));

	qlOBUF QL_INST_F2A_B_4_5 (.IN_OBUF(m1_oper0_wdata_dup_0[30]),.OUT_OBUF(m1_oper0_wdata[30]));

	qlOBUF QL_INST_F2A_B_4_6 (.IN_OBUF(m1_oper0_wdata_dup_0[29]),.OUT_OBUF(m1_oper0_wdata[29]));

	qlOBUF QL_INST_F2A_B_4_7 (.IN_OBUF(m1_oper0_wdata_dup_0[28]),.OUT_OBUF(m1_oper0_wdata[28]));

	qlOBUF QL_INST_F2A_B_4_8 (.IN_OBUF(m1_oper0_wdata_dup_0[27]),.OUT_OBUF(m1_oper0_wdata[27]));

	qlOBUF QL_INST_F2A_B_4_9 (.IN_OBUF(m1_oper0_wdata_dup_0[26]),.OUT_OBUF(m1_oper0_wdata[26]));

	qlOBUF QL_INST_F2A_B_4_10 (.IN_OBUF(m1_oper0_wdata_dup_0[25]),.OUT_OBUF(m1_oper0_wdata[25]));

	qlOBUF QL_INST_F2A_B_4_11 (.IN_OBUF(m1_oper0_wdata_dup_0[24]),.OUT_OBUF(m1_oper0_wdata[24]));

	qlOBUF QL_INST_F2A_B_4_12 (.IN_OBUF(m1_oper0_wdata_dup_0[23]),.OUT_OBUF(m1_oper0_wdata[23]));

	qlOBUF QL_INST_F2A_B_4_13 (.IN_OBUF(m1_oper0_wdata_dup_0[22]),.OUT_OBUF(m1_oper0_wdata[22]));

	qlOBUF QL_INST_F2A_B_4_14 (.IN_OBUF(m1_oper0_wdata_dup_0[21]),.OUT_OBUF(m1_oper0_wdata[21]));

	qlOBUF QL_INST_F2A_B_4_15 (.IN_OBUF(m1_oper0_wdata_dup_0[20]),.OUT_OBUF(m1_oper0_wdata[20]));

	qlOBUF QL_INST_F2A_B_4_16 (.IN_OBUF(m1_oper0_wdata_dup_0[19]),.OUT_OBUF(m1_oper0_wdata[19]));

	qlOBUF QL_INST_F2A_B_4_17 (.IN_OBUF(m1_oper0_wdata_dup_0[18]),.OUT_OBUF(m1_oper0_wdata[18]));

	qlIBUF QL_INST_A2F_B_4_0 (.IN_IBUF(m1_oper0_rdata[27]),.OUT_IBUF(m1_oper0_rdata_int[27]));

	qlIBUF QL_INST_A2F_B_4_1 (.IN_IBUF(m1_oper0_rdata[26]),.OUT_IBUF(m1_oper0_rdata_int[26]));

	qlIBUF QL_INST_A2F_B_4_2 (.IN_IBUF(m1_oper0_rdata[25]),.OUT_IBUF(m1_oper0_rdata_int[25]));

	qlIBUF QL_INST_A2F_B_4_3 (.IN_IBUF(m1_oper0_rdata[24]),.OUT_IBUF(m1_oper0_rdata_int[24]));

	qlIBUF QL_INST_A2F_B_4_4 (.IN_IBUF(m1_oper0_rdata[23]),.OUT_IBUF(m1_oper0_rdata_int[23]));

	qlIBUF QL_INST_A2F_B_4_5 (.IN_IBUF(m1_oper0_rdata[22]),.OUT_IBUF(m1_oper0_rdata_int[22]));

	qlIBUF QL_INST_A2F_B_4_6 (.IN_IBUF(m1_oper0_rdata[21]),.OUT_IBUF(m1_oper0_rdata_int[21]));

	qlIBUF QL_INST_A2F_B_4_7 (.IN_IBUF(m1_oper0_rdata[20]),.OUT_IBUF(m1_oper0_rdata_int[20]));

	qlOBUF QL_INST_F2A_B_5_0 (.IN_OBUF(m1_oper0_wdata_dup_0[17]),.OUT_OBUF(m1_oper0_wdata[17]));

	qlOBUF QL_INST_F2A_B_5_1 (.IN_OBUF(m1_oper0_wdata_dup_0[16]),.OUT_OBUF(m1_oper0_wdata[16]));

	qlOBUF QL_INST_F2A_B_5_2 (.IN_OBUF(m1_oper0_wdata_dup_0[15]),.OUT_OBUF(m1_oper0_wdata[15]));

	qlOBUF QL_INST_F2A_B_5_3 (.IN_OBUF(m1_oper0_wdata_dup_0[14]),.OUT_OBUF(m1_oper0_wdata[14]));

	qlOBUF QL_INST_F2A_B_5_4 (.IN_OBUF(m1_oper0_wdata_dup_0[13]),.OUT_OBUF(m1_oper0_wdata[13]));

	qlOBUF QL_INST_F2A_B_5_5 (.IN_OBUF(m1_oper0_wdata_dup_0[12]),.OUT_OBUF(m1_oper0_wdata[12]));

	qlOBUF QL_INST_F2A_B_5_6 (.IN_OBUF(m1_oper0_wdata_dup_0[11]),.OUT_OBUF(m1_oper0_wdata[11]));

	qlOBUF QL_INST_F2A_B_5_7 (.IN_OBUF(m1_oper0_wdata_dup_0[10]),.OUT_OBUF(m1_oper0_wdata[10]));

	qlOBUF QL_INST_F2A_B_5_8 (.IN_OBUF(m1_oper0_wdata_dup_0[9]),.OUT_OBUF(m1_oper0_wdata[9]));

	qlOBUF QL_INST_F2A_B_5_9 (.IN_OBUF(m1_oper0_wdata_dup_0[8]),.OUT_OBUF(m1_oper0_wdata[8]));

	qlOBUF QL_INST_F2A_B_5_10 (.IN_OBUF(m1_oper0_wdata_dup_0[7]),.OUT_OBUF(m1_oper0_wdata[7]));

	qlOBUF QL_INST_F2A_B_5_11 (.IN_OBUF(m1_oper0_wdata_dup_0[6]),.OUT_OBUF(m1_oper0_wdata[6]));

	qlIBUF QL_INST_A2F_B_5_0 (.IN_IBUF(m1_oper0_rdata[19]),.OUT_IBUF(m1_oper0_rdata_int[19]));

	qlIBUF QL_INST_A2F_B_5_1 (.IN_IBUF(m1_oper0_rdata[18]),.OUT_IBUF(m1_oper0_rdata_int[18]));

	qlIBUF QL_INST_A2F_B_5_2 (.IN_IBUF(m1_oper0_rdata[17]),.OUT_IBUF(m1_oper0_rdata_int[17]));

	qlIBUF QL_INST_A2F_B_5_3 (.IN_IBUF(m1_oper0_rdata[16]),.OUT_IBUF(m1_oper0_rdata_int[16]));

	qlIBUF QL_INST_A2F_B_5_4 (.IN_IBUF(m1_oper0_rdata[15]),.OUT_IBUF(m1_oper0_rdata_int[15]));

	qlIBUF QL_INST_A2F_B_5_5 (.IN_IBUF(m1_oper0_rdata[14]),.OUT_IBUF(m1_oper0_rdata_int[14]));

	qlOBUF QL_INST_F2A_B_6_0 (.IN_OBUF(m1_oper0_wdata_dup_0[5]),.OUT_OBUF(m1_oper0_wdata[5]));

	qlOBUF QL_INST_F2A_B_6_1 (.IN_OBUF(m1_oper0_wdata_dup_0[4]),.OUT_OBUF(m1_oper0_wdata[4]));

	qlOBUF QL_INST_F2A_B_6_2 (.IN_OBUF(m1_oper0_wdata_dup_0[3]),.OUT_OBUF(m1_oper0_wdata[3]));

	qlOBUF QL_INST_F2A_B_6_3 (.IN_OBUF(m1_oper0_wdata_dup_0[2]),.OUT_OBUF(m1_oper0_wdata[2]));

	qlOBUF QL_INST_F2A_B_6_4 (.IN_OBUF(m1_oper0_wdata_dup_0[1]),.OUT_OBUF(m1_oper0_wdata[1]));

	qlOBUF QL_INST_F2A_B_6_5 (.IN_OBUF(m1_oper0_wdata_dup_0[0]),.OUT_OBUF(m1_oper0_wdata[0]));

	qlOBUF QL_INST_F2A_B_6_7 (.IN_OBUF(m1_oper0_waddr_dup_0[11]),.OUT_OBUF(m1_oper0_waddr[11]));

	qlOBUF QL_INST_F2A_B_6_8 (.IN_OBUF(m1_oper0_waddr_dup_0[10]),.OUT_OBUF(m1_oper0_waddr[10]));

	qlOBUF QL_INST_F2A_B_6_9 (.IN_OBUF(m1_oper0_waddr_dup_0[9]),.OUT_OBUF(m1_oper0_waddr[9]));

	qlOBUF QL_INST_F2A_B_6_10 (.IN_OBUF(m1_oper0_waddr_dup_0[8]),.OUT_OBUF(m1_oper0_waddr[8]));

	qlOBUF QL_INST_F2A_B_6_11 (.IN_OBUF(m1_oper0_waddr_dup_0[7]),.OUT_OBUF(m1_oper0_waddr[7]));

	qlOBUF QL_INST_F2A_B_6_12 (.IN_OBUF(m1_oper0_waddr_dup_0[6]),.OUT_OBUF(m1_oper0_waddr[6]));

	qlOBUF QL_INST_F2A_B_6_13 (.IN_OBUF(m1_oper0_waddr_dup_0[5]),.OUT_OBUF(m1_oper0_waddr[5]));

	qlOBUF QL_INST_F2A_B_6_14 (.IN_OBUF(m1_oper0_waddr_dup_0[4]),.OUT_OBUF(m1_oper0_waddr[4]));

	qlOBUF QL_INST_F2A_B_6_15 (.IN_OBUF(m1_oper0_waddr_dup_0[3]),.OUT_OBUF(m1_oper0_waddr[3]));

	qlOBUF QL_INST_F2A_B_6_16 (.IN_OBUF(m1_oper0_waddr_dup_0[2]),.OUT_OBUF(m1_oper0_waddr[2]));

	qlOBUF QL_INST_F2A_B_6_17 (.IN_OBUF(m1_oper0_waddr_dup_0[1]),.OUT_OBUF(m1_oper0_waddr[1]));

	DBUF QL_INST_F2Adef_B_6_1 (.IN_DBUF(GND),.OUT_DBUF(m0_oper1_powerdn));

	qlIBUF QL_INST_A2F_B_6_0 (.IN_IBUF(m1_oper0_rdata[13]),.OUT_IBUF(m1_oper0_rdata_int[13]));

	qlIBUF QL_INST_A2F_B_6_1 (.IN_IBUF(m1_oper0_rdata[12]),.OUT_IBUF(m1_oper0_rdata_int[12]));

	qlIBUF QL_INST_A2F_B_6_2 (.IN_IBUF(m1_oper0_rdata[11]),.OUT_IBUF(m1_oper0_rdata_int[11]));

	qlIBUF QL_INST_A2F_B_6_3 (.IN_IBUF(m1_oper0_rdata[10]),.OUT_IBUF(m1_oper0_rdata_int[10]));

	qlIBUF QL_INST_A2F_B_6_4 (.IN_IBUF(m1_oper0_rdata[9]),.OUT_IBUF(m1_oper0_rdata_int[9]));

	qlIBUF QL_INST_A2F_B_6_5 (.IN_IBUF(m1_oper0_rdata[8]),.OUT_IBUF(m1_oper0_rdata_int[8]));

	qlIBUF QL_INST_A2F_B_6_6 (.IN_IBUF(m1_oper0_rdata[7]),.OUT_IBUF(m1_oper0_rdata_int[7]));

	qlIBUF QL_INST_A2F_B_6_7 (.IN_IBUF(m1_oper0_rdata[6]),.OUT_IBUF(m1_oper0_rdata_int[6]));

	qlOBUF QL_INST_F2A_B_7_0 (.IN_OBUF(m1_oper0_waddr_dup_0[0]),.OUT_OBUF(m1_oper0_waddr[0]));

	qlOBUF QL_INST_F2A_B_7_1 (.IN_OBUF(m1_oper0_we_dup_0),.OUT_OBUF(m1_oper0_we));

	qlOBUF QL_INST_F2A_B_7_2 (.IN_OBUF(m0_oper0_wdsel_dup_0),.OUT_OBUF(m1_oper0_wdsel));

	qlOBUF QL_INST_F2A_B_7_3 (.IN_OBUF(m0_oper0_rmode_dup_0[1]),.OUT_OBUF(m1_oper0_rmode[1]));

	qlOBUF QL_INST_F2A_B_7_4 (.IN_OBUF(m0_oper0_rmode_dup_0[0]),.OUT_OBUF(m1_oper0_rmode[0]));

	qlOBUF QL_INST_F2A_B_7_5 (.IN_OBUF(m1_oper0_raddr_dup_0[11]),.OUT_OBUF(m1_oper0_raddr[11]));

	qlOBUF QL_INST_F2A_B_7_6 (.IN_OBUF(m1_oper0_raddr_dup_0[10]),.OUT_OBUF(m1_oper0_raddr[10]));

	qlOBUF QL_INST_F2A_B_7_7 (.IN_OBUF(m1_oper0_raddr_dup_0[9]),.OUT_OBUF(m1_oper0_raddr[9]));

	qlOBUF QL_INST_F2A_B_7_8 (.IN_OBUF(m1_oper0_raddr_dup_0[8]),.OUT_OBUF(m1_oper0_raddr[8]));

	qlOBUF QL_INST_F2A_B_7_9 (.IN_OBUF(m1_oper0_raddr_dup_0[7]),.OUT_OBUF(m1_oper0_raddr[7]));

	qlOBUF QL_INST_F2A_B_7_10 (.IN_OBUF(m1_oper0_raddr_dup_0[6]),.OUT_OBUF(m1_oper0_raddr[6]));

	qlOBUF QL_INST_F2A_B_7_11 (.IN_OBUF(m1_oper0_raddr_dup_0[5]),.OUT_OBUF(m1_oper0_raddr[5]));

	qlIBUF QL_INST_A2F_B_7_0 (.IN_IBUF(m1_oper0_rdata[5]),.OUT_IBUF(m1_oper0_rdata_int[5]));

	qlIBUF QL_INST_A2F_B_7_1 (.IN_IBUF(m1_oper0_rdata[4]),.OUT_IBUF(m1_oper0_rdata_int[4]));

	qlIBUF QL_INST_A2F_B_7_2 (.IN_IBUF(m1_oper0_rdata[3]),.OUT_IBUF(m1_oper0_rdata_int[3]));

	qlIBUF QL_INST_A2F_B_7_3 (.IN_IBUF(m1_oper0_rdata[2]),.OUT_IBUF(m1_oper0_rdata_int[2]));

	qlIBUF QL_INST_A2F_B_7_4 (.IN_IBUF(m1_oper0_rdata[1]),.OUT_IBUF(m1_oper0_rdata_int[1]));

	qlIBUF QL_INST_A2F_B_7_5 (.IN_IBUF(m1_oper0_rdata[0]),.OUT_IBUF(m1_oper0_rdata_int[0]));

	qlOBUF QL_INST_F2A_B_8_0 (.IN_OBUF(CLK_int_0__CAND0_BLSBL_8_padClk),.OUT_OBUF(m1_oper0_rclk));

	qlOBUF QL_INST_F2A_B_8_1 (.IN_OBUF(m1_oper0_raddr_dup_0[4]),.OUT_OBUF(m1_oper0_raddr[4]));

	qlOBUF QL_INST_F2A_B_8_2 (.IN_OBUF(m1_oper0_raddr_dup_0[3]),.OUT_OBUF(m1_oper0_raddr[3]));

	qlOBUF QL_INST_F2A_B_8_3 (.IN_OBUF(m1_oper0_raddr_dup_0[2]),.OUT_OBUF(m1_oper0_raddr[2]));

	qlOBUF QL_INST_F2A_B_8_4 (.IN_OBUF(m1_oper0_raddr_dup_0[1]),.OUT_OBUF(m1_oper0_raddr[1]));

	qlOBUF QL_INST_F2A_B_8_5 (.IN_OBUF(m1_oper0_raddr_dup_0[0]),.OUT_OBUF(m1_oper0_raddr[0]));

	qlOBUF QL_INST_F2A_B_8_7 (.IN_OBUF(m1_m0_osel_dup_0),.OUT_OBUF(m1_m0_osel));

	qlOBUF QL_INST_F2A_B_8_8 (.IN_OBUF(m1_m0_clken_dup_0),.OUT_OBUF(m1_m0_clken));

	qlOBUF QL_INST_F2A_B_8_9 (.IN_OBUF(m1_m0_outsel_dup_0[5]),.OUT_OBUF(m1_m0_outsel[5]));

	qlOBUF QL_INST_F2A_B_8_10 (.IN_OBUF(m1_m0_outsel_dup_0[4]),.OUT_OBUF(m1_m0_outsel[4]));

	qlOBUF QL_INST_F2A_B_8_11 (.IN_OBUF(m1_m0_outsel_dup_0[3]),.OUT_OBUF(m1_m0_outsel[3]));

	qlOBUF QL_INST_F2A_B_8_12 (.IN_OBUF(m1_m0_outsel_dup_0[2]),.OUT_OBUF(m1_m0_outsel[2]));

	qlOBUF QL_INST_F2A_B_8_13 (.IN_OBUF(m1_m0_outsel_dup_0[1]),.OUT_OBUF(m1_m0_outsel[1]));

	qlOBUF QL_INST_F2A_B_8_14 (.IN_OBUF(m1_m0_outsel_dup_0[0]),.OUT_OBUF(m1_m0_outsel[0]));

	qlOBUF QL_INST_F2A_B_8_15 (.IN_OBUF(m1_m0_sat_dup_0),.OUT_OBUF(m1_m0_sat));

	qlOBUF QL_INST_F2A_B_8_16 (.IN_OBUF(m1_m0_rnd_dup_0),.OUT_OBUF(m1_m0_rnd));

	qlOBUF QL_INST_F2A_B_8_17 (.IN_OBUF(m1_m0_clr_dup_0),.OUT_OBUF(m1_m0_clr));

	qlIBUF QL_INST_A2F_B_8_4 (.IN_IBUF(m1_m0_dataout[31]),.OUT_IBUF(m1_m0_dataout_int[31]));

	qlIBUF QL_INST_A2F_B_8_5 (.IN_IBUF(m1_m0_dataout[30]),.OUT_IBUF(m1_m0_dataout_int[30]));

	qlIBUF QL_INST_A2F_B_8_6 (.IN_IBUF(m1_m0_dataout[29]),.OUT_IBUF(m1_m0_dataout_int[29]));

	qlIBUF QL_INST_A2F_B_8_7 (.IN_IBUF(m1_m0_dataout[28]),.OUT_IBUF(m1_m0_dataout_int[28]));

	qlOBUF QL_INST_F2A_B_9_0 (.IN_OBUF(CLK_int_0__CAND0_BLSBR_9_padClk),.OUT_OBUF(m1_m0_clk));

	qlOBUF QL_INST_F2A_B_9_1 (.IN_OBUF(m1_oper0_rdata_int[31]),.OUT_OBUF(m1_m0_oper_in[31]));

	qlOBUF QL_INST_F2A_B_9_2 (.IN_OBUF(m1_oper0_rdata_int[30]),.OUT_OBUF(m1_m0_oper_in[30]));

	qlOBUF QL_INST_F2A_B_9_3 (.IN_OBUF(m1_oper0_rdata_int[29]),.OUT_OBUF(m1_m0_oper_in[29]));

	qlOBUF QL_INST_F2A_B_9_4 (.IN_OBUF(m1_oper0_rdata_int[28]),.OUT_OBUF(m1_m0_oper_in[28]));

	qlOBUF QL_INST_F2A_B_9_5 (.IN_OBUF(m1_oper0_rdata_int[27]),.OUT_OBUF(m1_m0_oper_in[27]));

	qlOBUF QL_INST_F2A_B_9_6 (.IN_OBUF(m1_oper0_rdata_int[26]),.OUT_OBUF(m1_m0_oper_in[26]));

	qlOBUF QL_INST_F2A_B_9_7 (.IN_OBUF(m1_oper0_rdata_int[25]),.OUT_OBUF(m1_m0_oper_in[25]));

	qlOBUF QL_INST_F2A_B_9_8 (.IN_OBUF(m1_oper0_rdata_int[24]),.OUT_OBUF(m1_m0_oper_in[24]));

	qlOBUF QL_INST_F2A_B_9_9 (.IN_OBUF(m1_oper0_rdata_int[23]),.OUT_OBUF(m1_m0_oper_in[23]));

	qlOBUF QL_INST_F2A_B_9_10 (.IN_OBUF(m1_oper0_rdata_int[22]),.OUT_OBUF(m1_m0_oper_in[22]));

	qlOBUF QL_INST_F2A_B_9_11 (.IN_OBUF(m1_oper0_rdata_int[21]),.OUT_OBUF(m1_m0_oper_in[21]));

	qlIBUF QL_INST_A2F_B_9_0 (.IN_IBUF(m1_m0_dataout[27]),.OUT_IBUF(m1_m0_dataout_int[27]));

	qlIBUF QL_INST_A2F_B_9_1 (.IN_IBUF(m1_m0_dataout[26]),.OUT_IBUF(m1_m0_dataout_int[26]));

	qlIBUF QL_INST_A2F_B_9_2 (.IN_IBUF(m1_m0_dataout[25]),.OUT_IBUF(m1_m0_dataout_int[25]));

	qlIBUF QL_INST_A2F_B_9_3 (.IN_IBUF(m1_m0_dataout[24]),.OUT_IBUF(m1_m0_dataout_int[24]));

	qlIBUF QL_INST_A2F_B_9_4 (.IN_IBUF(m1_m0_dataout[23]),.OUT_IBUF(m1_m0_dataout_int[23]));

	qlIBUF QL_INST_A2F_B_9_5 (.IN_IBUF(m1_m0_dataout[22]),.OUT_IBUF(m1_m0_dataout_int[22]));

	qlOBUF QL_INST_F2A_B_10_0 (.IN_OBUF(m1_oper0_rdata_int[20]),.OUT_OBUF(m1_m0_oper_in[20]));

	qlOBUF QL_INST_F2A_B_10_1 (.IN_OBUF(m1_oper0_rdata_int[19]),.OUT_OBUF(m1_m0_oper_in[19]));

	qlOBUF QL_INST_F2A_B_10_2 (.IN_OBUF(m1_oper0_rdata_int[18]),.OUT_OBUF(m1_m0_oper_in[18]));

	qlOBUF QL_INST_F2A_B_10_3 (.IN_OBUF(m1_oper0_rdata_int[17]),.OUT_OBUF(m1_m0_oper_in[17]));

	qlOBUF QL_INST_F2A_B_10_4 (.IN_OBUF(m1_oper0_rdata_int[16]),.OUT_OBUF(m1_m0_oper_in[16]));

	qlOBUF QL_INST_F2A_B_10_5 (.IN_OBUF(m1_oper0_rdata_int[15]),.OUT_OBUF(m1_m0_oper_in[15]));

	qlOBUF QL_INST_F2A_B_10_6 (.IN_OBUF(m1_oper0_rdata_int[14]),.OUT_OBUF(m1_m0_oper_in[14]));

	qlOBUF QL_INST_F2A_B_10_7 (.IN_OBUF(m1_oper0_rdata_int[13]),.OUT_OBUF(m1_m0_oper_in[13]));

	qlOBUF QL_INST_F2A_B_10_8 (.IN_OBUF(m1_oper0_rdata_int[12]),.OUT_OBUF(m1_m0_oper_in[12]));

	qlOBUF QL_INST_F2A_B_10_9 (.IN_OBUF(m1_oper0_rdata_int[11]),.OUT_OBUF(m1_m0_oper_in[11]));

	qlOBUF QL_INST_F2A_B_10_10 (.IN_OBUF(m1_oper0_rdata_int[10]),.OUT_OBUF(m1_m0_oper_in[10]));

	qlOBUF QL_INST_F2A_B_10_11 (.IN_OBUF(m1_oper0_rdata_int[9]),.OUT_OBUF(m1_m0_oper_in[9]));

	qlOBUF QL_INST_F2A_B_10_12 (.IN_OBUF(m1_oper0_rdata_int[8]),.OUT_OBUF(m1_m0_oper_in[8]));

	qlOBUF QL_INST_F2A_B_10_13 (.IN_OBUF(m1_oper0_rdata_int[7]),.OUT_OBUF(m1_m0_oper_in[7]));

	qlOBUF QL_INST_F2A_B_10_14 (.IN_OBUF(m1_oper0_rdata_int[6]),.OUT_OBUF(m1_m0_oper_in[6]));

	qlOBUF QL_INST_F2A_B_10_15 (.IN_OBUF(m1_oper0_rdata_int[5]),.OUT_OBUF(m1_m0_oper_in[5]));

	qlOBUF QL_INST_F2A_B_10_16 (.IN_OBUF(m1_oper0_rdata_int[4]),.OUT_OBUF(m1_m0_oper_in[4]));

	qlOBUF QL_INST_F2A_B_10_17 (.IN_OBUF(m1_oper0_rdata_int[3]),.OUT_OBUF(m1_m0_oper_in[3]));

	qlIBUF QL_INST_A2F_B_10_0 (.IN_IBUF(m1_m0_dataout[21]),.OUT_IBUF(m1_m0_dataout_int[21]));

	qlIBUF QL_INST_A2F_B_10_1 (.IN_IBUF(m1_m0_dataout[20]),.OUT_IBUF(m1_m0_dataout_int[20]));

	qlIBUF QL_INST_A2F_B_10_2 (.IN_IBUF(m1_m0_dataout[19]),.OUT_IBUF(m1_m0_dataout_int[19]));

	qlIBUF QL_INST_A2F_B_10_3 (.IN_IBUF(m1_m0_dataout[18]),.OUT_IBUF(m1_m0_dataout_int[18]));

	qlIBUF QL_INST_A2F_B_10_4 (.IN_IBUF(m1_m0_dataout[17]),.OUT_IBUF(m1_m0_dataout_int[17]));

	qlIBUF QL_INST_A2F_B_10_5 (.IN_IBUF(m1_m0_dataout[16]),.OUT_IBUF(m1_m0_dataout_int[16]));

	qlIBUF QL_INST_A2F_B_10_6 (.IN_IBUF(m1_m0_dataout[15]),.OUT_IBUF(m1_m0_dataout_int[15]));

	qlIBUF QL_INST_A2F_B_10_7 (.IN_IBUF(m1_m0_dataout[14]),.OUT_IBUF(m1_m0_dataout_int[14]));

	qlOBUF QL_INST_F2A_B_11_0 (.IN_OBUF(m1_oper0_rdata_int[2]),.OUT_OBUF(m1_m0_oper_in[2]));

	qlOBUF QL_INST_F2A_B_11_1 (.IN_OBUF(m1_oper0_rdata_int[1]),.OUT_OBUF(m1_m0_oper_in[1]));

	qlOBUF QL_INST_F2A_B_11_2 (.IN_OBUF(m1_oper0_rdata_int[0]),.OUT_OBUF(m1_m0_oper_in[0]));

	qlOBUF QL_INST_F2A_B_11_3 (.IN_OBUF(m1_m0_csel_dup_0),.OUT_OBUF(m1_m0_csel));

	qlOBUF QL_INST_F2A_B_11_4 (.IN_OBUF(m1_coef_rdata_int[31]),.OUT_OBUF(m1_m0_coef_in[31]));

	qlOBUF QL_INST_F2A_B_11_5 (.IN_OBUF(m1_coef_rdata_int[30]),.OUT_OBUF(m1_m0_coef_in[30]));

	qlOBUF QL_INST_F2A_B_11_6 (.IN_OBUF(m1_coef_rdata_int[29]),.OUT_OBUF(m1_m0_coef_in[29]));

	qlOBUF QL_INST_F2A_B_11_7 (.IN_OBUF(m1_coef_rdata_int[28]),.OUT_OBUF(m1_m0_coef_in[28]));

	qlOBUF QL_INST_F2A_B_11_8 (.IN_OBUF(m1_coef_rdata_int[27]),.OUT_OBUF(m1_m0_coef_in[27]));

	qlOBUF QL_INST_F2A_B_11_9 (.IN_OBUF(m1_coef_rdata_int[26]),.OUT_OBUF(m1_m0_coef_in[26]));

	qlOBUF QL_INST_F2A_B_11_10 (.IN_OBUF(m1_coef_rdata_int[25]),.OUT_OBUF(m1_m0_coef_in[25]));

	qlOBUF QL_INST_F2A_B_11_11 (.IN_OBUF(m1_coef_rdata_int[24]),.OUT_OBUF(m1_m0_coef_in[24]));

	qlIBUF QL_INST_A2F_B_11_0 (.IN_IBUF(m1_m0_dataout[13]),.OUT_IBUF(m1_m0_dataout_int[13]));

	qlIBUF QL_INST_A2F_B_11_1 (.IN_IBUF(m1_m0_dataout[12]),.OUT_IBUF(m1_m0_dataout_int[12]));

	qlIBUF QL_INST_A2F_B_11_2 (.IN_IBUF(m1_m0_dataout[11]),.OUT_IBUF(m1_m0_dataout_int[11]));

	qlIBUF QL_INST_A2F_B_11_3 (.IN_IBUF(m1_m0_dataout[10]),.OUT_IBUF(m1_m0_dataout_int[10]));

	qlIBUF QL_INST_A2F_B_11_4 (.IN_IBUF(m1_m0_dataout[9]),.OUT_IBUF(m1_m0_dataout_int[9]));

	qlIBUF QL_INST_A2F_B_11_5 (.IN_IBUF(m1_m0_dataout[8]),.OUT_IBUF(m1_m0_dataout_int[8]));

	qlOBUF QL_INST_F2A_B_12_0 (.IN_OBUF(m1_coef_rdata_int[23]),.OUT_OBUF(m1_m0_coef_in[23]));

	qlOBUF QL_INST_F2A_B_12_1 (.IN_OBUF(m1_coef_rdata_int[22]),.OUT_OBUF(m1_m0_coef_in[22]));

	qlOBUF QL_INST_F2A_B_12_2 (.IN_OBUF(m1_coef_rdata_int[21]),.OUT_OBUF(m1_m0_coef_in[21]));

	qlOBUF QL_INST_F2A_B_12_3 (.IN_OBUF(m1_coef_rdata_int[20]),.OUT_OBUF(m1_m0_coef_in[20]));

	qlOBUF QL_INST_F2A_B_12_4 (.IN_OBUF(m1_coef_rdata_int[19]),.OUT_OBUF(m1_m0_coef_in[19]));

	qlOBUF QL_INST_F2A_B_12_5 (.IN_OBUF(m1_coef_rdata_int[18]),.OUT_OBUF(m1_m0_coef_in[18]));

	qlOBUF QL_INST_F2A_B_12_6 (.IN_OBUF(m1_coef_rdata_int[17]),.OUT_OBUF(m1_m0_coef_in[17]));

	qlOBUF QL_INST_F2A_B_12_7 (.IN_OBUF(m1_coef_rdata_int[16]),.OUT_OBUF(m1_m0_coef_in[16]));

	qlOBUF QL_INST_F2A_B_12_8 (.IN_OBUF(m1_coef_rdata_int[15]),.OUT_OBUF(m1_m0_coef_in[15]));

	qlOBUF QL_INST_F2A_B_12_9 (.IN_OBUF(m1_coef_rdata_int[14]),.OUT_OBUF(m1_m0_coef_in[14]));

	qlOBUF QL_INST_F2A_B_12_10 (.IN_OBUF(m1_coef_rdata_int[13]),.OUT_OBUF(m1_m0_coef_in[13]));

	qlOBUF QL_INST_F2A_B_12_11 (.IN_OBUF(m1_coef_rdata_int[12]),.OUT_OBUF(m1_m0_coef_in[12]));

	qlOBUF QL_INST_F2A_B_12_12 (.IN_OBUF(m1_coef_rdata_int[11]),.OUT_OBUF(m1_m0_coef_in[11]));

	qlOBUF QL_INST_F2A_B_12_13 (.IN_OBUF(m1_coef_rdata_int[10]),.OUT_OBUF(m1_m0_coef_in[10]));

	qlOBUF QL_INST_F2A_B_12_14 (.IN_OBUF(m1_coef_rdata_int[9]),.OUT_OBUF(m1_m0_coef_in[9]));

	qlOBUF QL_INST_F2A_B_12_15 (.IN_OBUF(m1_coef_rdata_int[8]),.OUT_OBUF(m1_m0_coef_in[8]));

	qlOBUF QL_INST_F2A_B_12_16 (.IN_OBUF(m1_coef_rdata_int[7]),.OUT_OBUF(m1_m0_coef_in[7]));

	qlOBUF QL_INST_F2A_B_12_17 (.IN_OBUF(m1_coef_rdata_int[6]),.OUT_OBUF(m1_m0_coef_in[6]));

	qlIBUF QL_INST_A2F_B_12_0 (.IN_IBUF(m1_m0_dataout[7]),.OUT_IBUF(m1_m0_dataout_int[7]));

	qlIBUF QL_INST_A2F_B_12_1 (.IN_IBUF(m1_m0_dataout[6]),.OUT_IBUF(m1_m0_dataout_int[6]));

	qlIBUF QL_INST_A2F_B_12_2 (.IN_IBUF(m1_m0_dataout[5]),.OUT_IBUF(m1_m0_dataout_int[5]));

	qlIBUF QL_INST_A2F_B_12_3 (.IN_IBUF(m1_m0_dataout[4]),.OUT_IBUF(m1_m0_dataout_int[4]));

	qlIBUF QL_INST_A2F_B_12_4 (.IN_IBUF(m1_m0_dataout[3]),.OUT_IBUF(m1_m0_dataout_int[3]));

	qlIBUF QL_INST_A2F_B_12_5 (.IN_IBUF(m1_m0_dataout[2]),.OUT_IBUF(m1_m0_dataout_int[2]));

	qlIBUF QL_INST_A2F_B_12_6 (.IN_IBUF(m1_m0_dataout[1]),.OUT_IBUF(m1_m0_dataout_int[1]));

	qlIBUF QL_INST_A2F_B_12_7 (.IN_IBUF(m1_m0_dataout[0]),.OUT_IBUF(m1_m0_dataout_int[0]));

	qlOBUF QL_INST_F2A_B_13_0 (.IN_OBUF(m1_coef_rdata_int[5]),.OUT_OBUF(m1_m0_coef_in[5]));

	qlOBUF QL_INST_F2A_B_13_1 (.IN_OBUF(m1_coef_rdata_int[4]),.OUT_OBUF(m1_m0_coef_in[4]));

	qlOBUF QL_INST_F2A_B_13_2 (.IN_OBUF(m1_coef_rdata_int[3]),.OUT_OBUF(m1_m0_coef_in[3]));

	qlOBUF QL_INST_F2A_B_13_3 (.IN_OBUF(m1_coef_rdata_int[2]),.OUT_OBUF(m1_m0_coef_in[2]));

	qlOBUF QL_INST_F2A_B_13_4 (.IN_OBUF(m1_coef_rdata_int[1]),.OUT_OBUF(m1_m0_coef_in[1]));

	qlOBUF QL_INST_F2A_B_13_5 (.IN_OBUF(m1_coef_rdata_int[0]),.OUT_OBUF(m1_m0_coef_in[0]));

	qlOBUF QL_INST_F2A_B_13_6 (.IN_OBUF(m1_m0_mode_dup_0[1]),.OUT_OBUF(m1_m0_mode[1]));

	qlOBUF QL_INST_F2A_B_13_7 (.IN_OBUF(m1_m0_mode_dup_0[0]),.OUT_OBUF(m1_m0_mode[0]));

	qlOBUF QL_INST_F2A_B_13_8 (.IN_OBUF(m1_m0_tc_dup_0),.OUT_OBUF(m1_m0_tc));

	qlOBUF QL_INST_F2A_B_13_9 (.IN_OBUF(m1_m0_reset_dup_0),.OUT_OBUF(m1_m0_reset));

	qlOBUF QL_INST_F2A_B_13_10 (.IN_OBUF(m1_coef_wdata_dup_0[31]),.OUT_OBUF(m1_coef_wdata[31]));

	qlOBUF QL_INST_F2A_B_13_11 (.IN_OBUF(m1_coef_wdata_dup_0[30]),.OUT_OBUF(m1_coef_wdata[30]));

	qlIBUF QL_INST_A2F_B_13_2 (.IN_IBUF(m1_coef_rdata[31]),.OUT_IBUF(m1_coef_rdata_int[31]));

	qlIBUF QL_INST_A2F_B_13_3 (.IN_IBUF(m1_coef_rdata[30]),.OUT_IBUF(m1_coef_rdata_int[30]));

	qlIBUF QL_INST_A2F_B_13_4 (.IN_IBUF(m1_coef_rdata[29]),.OUT_IBUF(m1_coef_rdata_int[29]));

	qlIBUF QL_INST_A2F_B_13_5 (.IN_IBUF(m1_coef_rdata[28]),.OUT_IBUF(m1_coef_rdata_int[28]));

	qlOBUF QL_INST_F2A_B_14_0 (.IN_OBUF(m1_coef_wdata_dup_0[29]),.OUT_OBUF(m1_coef_wdata[29]));

	qlOBUF QL_INST_F2A_B_14_1 (.IN_OBUF(m1_coef_wdata_dup_0[28]),.OUT_OBUF(m1_coef_wdata[28]));

	qlOBUF QL_INST_F2A_B_14_2 (.IN_OBUF(m1_coef_wdata_dup_0[27]),.OUT_OBUF(m1_coef_wdata[27]));

	qlOBUF QL_INST_F2A_B_14_3 (.IN_OBUF(m1_coef_wdata_dup_0[26]),.OUT_OBUF(m1_coef_wdata[26]));

	qlOBUF QL_INST_F2A_B_14_4 (.IN_OBUF(m1_coef_wdata_dup_0[25]),.OUT_OBUF(m1_coef_wdata[25]));

	qlOBUF QL_INST_F2A_B_14_5 (.IN_OBUF(m1_coef_wdata_dup_0[24]),.OUT_OBUF(m1_coef_wdata[24]));

	qlOBUF QL_INST_F2A_B_14_6 (.IN_OBUF(m1_coef_wdata_dup_0[23]),.OUT_OBUF(m1_coef_wdata[23]));

	qlOBUF QL_INST_F2A_B_14_7 (.IN_OBUF(m1_coef_wdata_dup_0[22]),.OUT_OBUF(m1_coef_wdata[22]));

	qlOBUF QL_INST_F2A_B_14_8 (.IN_OBUF(m1_coef_wdata_dup_0[21]),.OUT_OBUF(m1_coef_wdata[21]));

	qlOBUF QL_INST_F2A_B_14_9 (.IN_OBUF(m1_coef_wdata_dup_0[20]),.OUT_OBUF(m1_coef_wdata[20]));

	qlOBUF QL_INST_F2A_B_14_10 (.IN_OBUF(m1_coef_wdata_dup_0[19]),.OUT_OBUF(m1_coef_wdata[19]));

	qlOBUF QL_INST_F2A_B_14_11 (.IN_OBUF(m1_coef_wdata_dup_0[18]),.OUT_OBUF(m1_coef_wdata[18]));

	qlOBUF QL_INST_F2A_B_14_12 (.IN_OBUF(m1_coef_wdata_dup_0[17]),.OUT_OBUF(m1_coef_wdata[17]));

	qlOBUF QL_INST_F2A_B_14_13 (.IN_OBUF(m1_coef_wdata_dup_0[16]),.OUT_OBUF(m1_coef_wdata[16]));

	qlOBUF QL_INST_F2A_B_14_14 (.IN_OBUF(m1_coef_wdata_dup_0[15]),.OUT_OBUF(m1_coef_wdata[15]));

	qlOBUF QL_INST_F2A_B_14_15 (.IN_OBUF(m1_coef_wdata_dup_0[14]),.OUT_OBUF(m1_coef_wdata[14]));

	qlOBUF QL_INST_F2A_B_14_16 (.IN_OBUF(m1_coef_wdata_dup_0[13]),.OUT_OBUF(m1_coef_wdata[13]));

	qlOBUF QL_INST_F2A_B_14_17 (.IN_OBUF(m1_coef_wdata_dup_0[12]),.OUT_OBUF(m1_coef_wdata[12]));

	qlIBUF QL_INST_A2F_B_14_0 (.IN_IBUF(m1_coef_rdata[27]),.OUT_IBUF(m1_coef_rdata_int[27]));

	qlIBUF QL_INST_A2F_B_14_1 (.IN_IBUF(m1_coef_rdata[26]),.OUT_IBUF(m1_coef_rdata_int[26]));

	qlIBUF QL_INST_A2F_B_14_2 (.IN_IBUF(m1_coef_rdata[25]),.OUT_IBUF(m1_coef_rdata_int[25]));

	qlIBUF QL_INST_A2F_B_14_3 (.IN_IBUF(m1_coef_rdata[24]),.OUT_IBUF(m1_coef_rdata_int[24]));

	qlIBUF QL_INST_A2F_B_14_4 (.IN_IBUF(m1_coef_rdata[23]),.OUT_IBUF(m1_coef_rdata_int[23]));

	qlIBUF QL_INST_A2F_B_14_5 (.IN_IBUF(m1_coef_rdata[22]),.OUT_IBUF(m1_coef_rdata_int[22]));

	qlIBUF QL_INST_A2F_B_14_6 (.IN_IBUF(m1_coef_rdata[21]),.OUT_IBUF(m1_coef_rdata_int[21]));

	qlIBUF QL_INST_A2F_B_14_7 (.IN_IBUF(m1_coef_rdata[20]),.OUT_IBUF(m1_coef_rdata_int[20]));

	qlOBUF QL_INST_F2A_B_15_0 (.IN_OBUF(m1_coef_wdata_dup_0[11]),.OUT_OBUF(m1_coef_wdata[11]));

	qlOBUF QL_INST_F2A_B_15_1 (.IN_OBUF(m1_coef_wdata_dup_0[10]),.OUT_OBUF(m1_coef_wdata[10]));

	qlOBUF QL_INST_F2A_B_15_2 (.IN_OBUF(m1_coef_wdata_dup_0[9]),.OUT_OBUF(m1_coef_wdata[9]));

	qlOBUF QL_INST_F2A_B_15_3 (.IN_OBUF(m1_coef_wdata_dup_0[8]),.OUT_OBUF(m1_coef_wdata[8]));

	qlOBUF QL_INST_F2A_B_15_4 (.IN_OBUF(m1_coef_wdata_dup_0[7]),.OUT_OBUF(m1_coef_wdata[7]));

	qlOBUF QL_INST_F2A_B_15_5 (.IN_OBUF(m1_coef_wdata_dup_0[6]),.OUT_OBUF(m1_coef_wdata[6]));

	qlOBUF QL_INST_F2A_B_15_6 (.IN_OBUF(m1_coef_wdata_dup_0[5]),.OUT_OBUF(m1_coef_wdata[5]));

	qlOBUF QL_INST_F2A_B_15_7 (.IN_OBUF(m1_coef_wdata_dup_0[4]),.OUT_OBUF(m1_coef_wdata[4]));

	qlOBUF QL_INST_F2A_B_15_8 (.IN_OBUF(m1_coef_wdata_dup_0[3]),.OUT_OBUF(m1_coef_wdata[3]));

	qlOBUF QL_INST_F2A_B_15_9 (.IN_OBUF(m1_coef_wdata_dup_0[2]),.OUT_OBUF(m1_coef_wdata[2]));

	qlOBUF QL_INST_F2A_B_15_10 (.IN_OBUF(m1_coef_wdata_dup_0[1]),.OUT_OBUF(m1_coef_wdata[1]));

	qlOBUF QL_INST_F2A_B_15_11 (.IN_OBUF(m1_coef_wdata_dup_0[0]),.OUT_OBUF(m1_coef_wdata[0]));

	qlIBUF QL_INST_A2F_B_15_0 (.IN_IBUF(m1_coef_rdata[19]),.OUT_IBUF(m1_coef_rdata_int[19]));

	qlIBUF QL_INST_A2F_B_15_1 (.IN_IBUF(m1_coef_rdata[18]),.OUT_IBUF(m1_coef_rdata_int[18]));

	qlIBUF QL_INST_A2F_B_15_2 (.IN_IBUF(m1_coef_rdata[17]),.OUT_IBUF(m1_coef_rdata_int[17]));

	qlIBUF QL_INST_A2F_B_15_3 (.IN_IBUF(m1_coef_rdata[16]),.OUT_IBUF(m1_coef_rdata_int[16]));

	qlIBUF QL_INST_A2F_B_15_4 (.IN_IBUF(m1_coef_rdata[15]),.OUT_IBUF(m1_coef_rdata_int[15]));

	qlIBUF QL_INST_A2F_B_15_5 (.IN_IBUF(m1_coef_rdata[14]),.OUT_IBUF(m1_coef_rdata_int[14]));

	qlOBUF QL_INST_F2A_B_16_0 (.IN_OBUF(CLK_int_0__CAND0_BLSBR_16_padClk),.OUT_OBUF(m1_coef_wclk));

	qlOBUF QL_INST_F2A_B_16_1 (.IN_OBUF(m1_coef_waddr_dup_0[11]),.OUT_OBUF(m1_coef_waddr[11]));

	qlOBUF QL_INST_F2A_B_16_2 (.IN_OBUF(m1_coef_waddr_dup_0[10]),.OUT_OBUF(m1_coef_waddr[10]));

	qlOBUF QL_INST_F2A_B_16_3 (.IN_OBUF(m1_coef_waddr_dup_0[9]),.OUT_OBUF(m1_coef_waddr[9]));

	qlOBUF QL_INST_F2A_B_16_4 (.IN_OBUF(m1_coef_waddr_dup_0[8]),.OUT_OBUF(m1_coef_waddr[8]));

	qlOBUF QL_INST_F2A_B_16_5 (.IN_OBUF(m1_coef_waddr_dup_0[7]),.OUT_OBUF(m1_coef_waddr[7]));

	qlOBUF QL_INST_F2A_B_16_6 (.IN_OBUF(m1_coef_waddr_dup_0[6]),.OUT_OBUF(m1_coef_waddr[6]));

	qlOBUF QL_INST_F2A_B_16_7 (.IN_OBUF(m1_coef_waddr_dup_0[5]),.OUT_OBUF(m1_coef_waddr[5]));

	qlOBUF QL_INST_F2A_B_16_8 (.IN_OBUF(m1_coef_waddr_dup_0[4]),.OUT_OBUF(m1_coef_waddr[4]));

	qlOBUF QL_INST_F2A_B_16_9 (.IN_OBUF(m1_coef_waddr_dup_0[3]),.OUT_OBUF(m1_coef_waddr[3]));

	qlOBUF QL_INST_F2A_B_16_10 (.IN_OBUF(m1_coef_waddr_dup_0[2]),.OUT_OBUF(m1_coef_waddr[2]));

	qlOBUF QL_INST_F2A_B_16_11 (.IN_OBUF(m1_coef_waddr_dup_0[1]),.OUT_OBUF(m1_coef_waddr[1]));

	qlOBUF QL_INST_F2A_B_16_12 (.IN_OBUF(m1_coef_waddr_dup_0[0]),.OUT_OBUF(m1_coef_waddr[0]));

	qlOBUF QL_INST_F2A_B_16_13 (.IN_OBUF(m1_coef_we_dup_0),.OUT_OBUF(m1_coef_we));

	qlIBUF QL_INST_A2F_B_16_3 (.IN_IBUF(m1_coef_rdata[13]),.OUT_IBUF(m1_coef_rdata_int[13]));

	qlIBUF QL_INST_A2F_B_16_4 (.IN_IBUF(m1_coef_rdata[12]),.OUT_IBUF(m1_coef_rdata_int[12]));

	qlIBUF QL_INST_A2F_B_16_5 (.IN_IBUF(m1_coef_rdata[11]),.OUT_IBUF(m1_coef_rdata_int[11]));

	qlIBUF QL_INST_A2F_B_16_6 (.IN_IBUF(m1_coef_rdata[10]),.OUT_IBUF(m1_coef_rdata_int[10]));

	qlIBUF QL_INST_A2F_B_16_7 (.IN_IBUF(m1_coef_rdata[9]),.OUT_IBUF(m1_coef_rdata_int[9]));

	qlOBUF QL_INST_F2A_B_17_0 (.IN_OBUF(CLK_int_0__CAND0_BRSBL_17_padClk),.OUT_OBUF(m1_coef_rclk));

	qlOBUF QL_INST_F2A_B_17_1 (.IN_OBUF(m1_coef_raddr_dup_0[11]),.OUT_OBUF(m1_coef_raddr[11]));

	qlOBUF QL_INST_F2A_B_17_2 (.IN_OBUF(m1_coef_raddr_dup_0[10]),.OUT_OBUF(m1_coef_raddr[10]));

	qlOBUF QL_INST_F2A_B_17_3 (.IN_OBUF(m1_coef_raddr_dup_0[9]),.OUT_OBUF(m1_coef_raddr[9]));

	qlOBUF QL_INST_F2A_B_17_4 (.IN_OBUF(m1_coef_raddr_dup_0[8]),.OUT_OBUF(m1_coef_raddr[8]));

	qlOBUF QL_INST_F2A_B_17_5 (.IN_OBUF(m1_coef_raddr_dup_0[7]),.OUT_OBUF(m1_coef_raddr[7]));

	qlOBUF QL_INST_F2A_B_17_6 (.IN_OBUF(m1_coef_raddr_dup_0[6]),.OUT_OBUF(m1_coef_raddr[6]));

	qlOBUF QL_INST_F2A_B_17_7 (.IN_OBUF(m1_coef_raddr_dup_0[5]),.OUT_OBUF(m1_coef_raddr[5]));

	qlOBUF QL_INST_F2A_B_17_8 (.IN_OBUF(m1_coef_raddr_dup_0[4]),.OUT_OBUF(m1_coef_raddr[4]));

	qlOBUF QL_INST_F2A_B_17_9 (.IN_OBUF(m0_coef_wdsel_dup_0),.OUT_OBUF(m1_coef_wdsel));

	qlOBUF QL_INST_F2A_B_17_10 (.IN_OBUF(m0_coef_rmode_dup_0[1]),.OUT_OBUF(m1_coef_rmode[1]));

	qlOBUF QL_INST_F2A_B_17_11 (.IN_OBUF(m0_coef_rmode_dup_0[0]),.OUT_OBUF(m1_coef_rmode[0]));

	qlIBUF QL_INST_A2F_B_17_0 (.IN_IBUF(m1_coef_rdata[5]),.OUT_IBUF(m1_coef_rdata_int[5]));

	qlIBUF QL_INST_A2F_B_17_1 (.IN_IBUF(m1_coef_rdata[4]),.OUT_IBUF(m1_coef_rdata_int[4]));

	qlIBUF QL_INST_A2F_B_17_2 (.IN_IBUF(m1_coef_rdata[3]),.OUT_IBUF(m1_coef_rdata_int[3]));

	qlIBUF QL_INST_A2F_B_17_3 (.IN_IBUF(m1_coef_rdata[8]),.OUT_IBUF(m1_coef_rdata_int[8]));

	qlIBUF QL_INST_A2F_B_17_4 (.IN_IBUF(m1_coef_rdata[7]),.OUT_IBUF(m1_coef_rdata_int[7]));

	qlIBUF QL_INST_A2F_B_17_5 (.IN_IBUF(m1_coef_rdata[6]),.OUT_IBUF(m1_coef_rdata_int[6]));

	qlOBUF QL_INST_F2A_B_18_0 (.IN_OBUF(m1_coef_raddr_dup_0[3]),.OUT_OBUF(m1_coef_raddr[3]));

	qlOBUF QL_INST_F2A_B_18_1 (.IN_OBUF(m1_coef_raddr_dup_0[2]),.OUT_OBUF(m1_coef_raddr[2]));

	qlOBUF QL_INST_F2A_B_18_2 (.IN_OBUF(m1_coef_raddr_dup_0[1]),.OUT_OBUF(m1_coef_raddr[1]));

	qlOBUF QL_INST_F2A_B_18_3 (.IN_OBUF(m1_coef_raddr_dup_0[0]),.OUT_OBUF(m1_coef_raddr[0]));

	qlOBUF QL_INST_F2A_B_18_4 (.IN_OBUF(m0_coef_wmode_dup_0[1]),.OUT_OBUF(m1_coef_wmode[1]));

	qlOBUF QL_INST_F2A_B_18_5 (.IN_OBUF(m0_coef_wmode_dup_0[0]),.OUT_OBUF(m1_coef_wmode[0]));

	qlOBUF QL_INST_F2A_B_18_7 (.IN_OBUF(m0_m0_outsel_dup_0[5]),.OUT_OBUF(m1_m1_outsel[5]));

	qlOBUF QL_INST_F2A_B_18_8 (.IN_OBUF(m0_m0_outsel_dup_0[4]),.OUT_OBUF(m1_m1_outsel[4]));

	qlOBUF QL_INST_F2A_B_18_9 (.IN_OBUF(m0_m0_outsel_dup_0[3]),.OUT_OBUF(m1_m1_outsel[3]));

	qlOBUF QL_INST_F2A_B_18_10 (.IN_OBUF(m0_m0_outsel_dup_0[2]),.OUT_OBUF(m1_m1_outsel[2]));

	qlOBUF QL_INST_F2A_B_18_11 (.IN_OBUF(m0_m0_outsel_dup_0[1]),.OUT_OBUF(m1_m1_outsel[1]));

	qlOBUF QL_INST_F2A_B_18_12 (.IN_OBUF(m0_m0_outsel_dup_0[0]),.OUT_OBUF(m1_m1_outsel[0]));

	qlOBUF QL_INST_F2A_B_18_13 (.IN_OBUF(m1_m1_sat_dup_0),.OUT_OBUF(m1_m1_sat));

	qlOBUF QL_INST_F2A_B_18_14 (.IN_OBUF(m1_m1_rnd_dup_0),.OUT_OBUF(m1_m1_rnd));

	qlOBUF QL_INST_F2A_B_18_15 (.IN_OBUF(m1_m1_clr_dup_0),.OUT_OBUF(m1_m1_clr));

	qlOBUF QL_INST_F2A_B_18_16 (.IN_OBUF(m1_m1_clken_dup_0),.OUT_OBUF(m1_m1_clken));

	DBUF QL_INST_F2Adef_B_18_1 (.IN_DBUF(GND),.OUT_DBUF(m0_coef_powerdn));

	qlIBUF QL_INST_A2F_B_18_0 (.IN_IBUF(m1_coef_rdata[2]),.OUT_IBUF(m1_coef_rdata_int[2]));

	qlIBUF QL_INST_A2F_B_18_1 (.IN_IBUF(m1_coef_rdata[1]),.OUT_IBUF(m1_coef_rdata_int[1]));

	qlIBUF QL_INST_A2F_B_18_2 (.IN_IBUF(m1_coef_rdata[0]),.OUT_IBUF(m1_coef_rdata_int[0]));

	qlIBUF QL_INST_A2F_B_18_6 (.IN_IBUF(m1_m1_dataout[31]),.OUT_IBUF(m1_m1_dataout_int[31]));

	qlIBUF QL_INST_A2F_B_18_7 (.IN_IBUF(m1_m1_dataout[30]),.OUT_IBUF(m1_m1_dataout_int[30]));

	qlOBUF QL_INST_F2A_B_19_0 (.IN_OBUF(CLK_int_0__CAND0_BRSBL_19_padClk),.OUT_OBUF(m1_m1_clk));

	qlOBUF QL_INST_F2A_B_19_1 (.IN_OBUF(m1_m1_osel_dup_0),.OUT_OBUF(m1_m1_osel));

	qlOBUF QL_INST_F2A_B_19_2 (.IN_OBUF(m1_m1_tc_dup_0),.OUT_OBUF(m1_m1_tc));

	qlOBUF QL_INST_F2A_B_19_3 (.IN_OBUF(m1_m1_reset_dup_0),.OUT_OBUF(m1_m1_reset));

	qlOBUF QL_INST_F2A_B_19_4 (.IN_OBUF(m1_coef_rdata_int[31]),.OUT_OBUF(m1_m1_coef_in[31]));

	qlOBUF QL_INST_F2A_B_19_5 (.IN_OBUF(m1_coef_rdata_int[30]),.OUT_OBUF(m1_m1_coef_in[30]));

	qlOBUF QL_INST_F2A_B_19_6 (.IN_OBUF(m1_coef_rdata_int[29]),.OUT_OBUF(m1_m1_coef_in[29]));

	qlOBUF QL_INST_F2A_B_19_7 (.IN_OBUF(m1_coef_rdata_int[28]),.OUT_OBUF(m1_m1_coef_in[28]));

	qlOBUF QL_INST_F2A_B_19_8 (.IN_OBUF(m1_coef_rdata_int[27]),.OUT_OBUF(m1_m1_coef_in[27]));

	qlOBUF QL_INST_F2A_B_19_9 (.IN_OBUF(m1_coef_rdata_int[26]),.OUT_OBUF(m1_m1_coef_in[26]));

	qlOBUF QL_INST_F2A_B_19_10 (.IN_OBUF(m1_coef_rdata_int[25]),.OUT_OBUF(m1_m1_coef_in[25]));

	qlOBUF QL_INST_F2A_B_19_11 (.IN_OBUF(m1_coef_rdata_int[24]),.OUT_OBUF(m1_m1_coef_in[24]));

	qlIBUF QL_INST_A2F_B_19_0 (.IN_IBUF(m1_m1_dataout[29]),.OUT_IBUF(m1_m1_dataout_int[29]));

	qlIBUF QL_INST_A2F_B_19_1 (.IN_IBUF(m1_m1_dataout[28]),.OUT_IBUF(m1_m1_dataout_int[28]));

	qlIBUF QL_INST_A2F_B_19_2 (.IN_IBUF(m1_m1_dataout[27]),.OUT_IBUF(m1_m1_dataout_int[27]));

	qlIBUF QL_INST_A2F_B_19_3 (.IN_IBUF(m1_m1_dataout[26]),.OUT_IBUF(m1_m1_dataout_int[26]));

	qlIBUF QL_INST_A2F_B_19_4 (.IN_IBUF(m1_m1_dataout[25]),.OUT_IBUF(m1_m1_dataout_int[25]));

	qlIBUF QL_INST_A2F_B_19_5 (.IN_IBUF(m1_m1_dataout[24]),.OUT_IBUF(m1_m1_dataout_int[24]));

	qlOBUF QL_INST_F2A_B_20_0 (.IN_OBUF(m1_coef_rdata_int[23]),.OUT_OBUF(m1_m1_coef_in[23]));

	qlOBUF QL_INST_F2A_B_20_1 (.IN_OBUF(m1_coef_rdata_int[22]),.OUT_OBUF(m1_m1_coef_in[22]));

	qlOBUF QL_INST_F2A_B_20_2 (.IN_OBUF(m1_coef_rdata_int[21]),.OUT_OBUF(m1_m1_coef_in[21]));

	qlOBUF QL_INST_F2A_B_20_3 (.IN_OBUF(m1_coef_rdata_int[20]),.OUT_OBUF(m1_m1_coef_in[20]));

	qlOBUF QL_INST_F2A_B_20_4 (.IN_OBUF(m1_coef_rdata_int[19]),.OUT_OBUF(m1_m1_coef_in[19]));

	qlOBUF QL_INST_F2A_B_20_5 (.IN_OBUF(m1_coef_rdata_int[18]),.OUT_OBUF(m1_m1_coef_in[18]));

	qlOBUF QL_INST_F2A_B_20_6 (.IN_OBUF(m1_coef_rdata_int[17]),.OUT_OBUF(m1_m1_coef_in[17]));

	qlOBUF QL_INST_F2A_B_20_7 (.IN_OBUF(m1_coef_rdata_int[16]),.OUT_OBUF(m1_m1_coef_in[16]));

	qlOBUF QL_INST_F2A_B_20_8 (.IN_OBUF(m1_coef_rdata_int[15]),.OUT_OBUF(m1_m1_coef_in[15]));

	qlOBUF QL_INST_F2A_B_20_9 (.IN_OBUF(m1_coef_rdata_int[14]),.OUT_OBUF(m1_m1_coef_in[14]));

	qlOBUF QL_INST_F2A_B_20_10 (.IN_OBUF(m1_coef_rdata_int[13]),.OUT_OBUF(m1_m1_coef_in[13]));

	qlOBUF QL_INST_F2A_B_20_11 (.IN_OBUF(m1_coef_rdata_int[12]),.OUT_OBUF(m1_m1_coef_in[12]));

	qlOBUF QL_INST_F2A_B_20_12 (.IN_OBUF(m1_coef_rdata_int[11]),.OUT_OBUF(m1_m1_coef_in[11]));

	qlOBUF QL_INST_F2A_B_20_13 (.IN_OBUF(m1_coef_rdata_int[10]),.OUT_OBUF(m1_m1_coef_in[10]));

	qlOBUF QL_INST_F2A_B_20_14 (.IN_OBUF(m1_coef_rdata_int[9]),.OUT_OBUF(m1_m1_coef_in[9]));

	qlOBUF QL_INST_F2A_B_20_15 (.IN_OBUF(m1_coef_rdata_int[8]),.OUT_OBUF(m1_m1_coef_in[8]));

	qlOBUF QL_INST_F2A_B_20_16 (.IN_OBUF(m1_coef_rdata_int[7]),.OUT_OBUF(m1_m1_coef_in[7]));

	qlOBUF QL_INST_F2A_B_20_17 (.IN_OBUF(m1_coef_rdata_int[6]),.OUT_OBUF(m1_m1_coef_in[6]));

	qlIBUF QL_INST_A2F_B_20_0 (.IN_IBUF(m1_m1_dataout[23]),.OUT_IBUF(m1_m1_dataout_int[23]));

	qlIBUF QL_INST_A2F_B_20_1 (.IN_IBUF(m1_m1_dataout[22]),.OUT_IBUF(m1_m1_dataout_int[22]));

	qlIBUF QL_INST_A2F_B_20_2 (.IN_IBUF(m1_m1_dataout[21]),.OUT_IBUF(m1_m1_dataout_int[21]));

	qlIBUF QL_INST_A2F_B_20_3 (.IN_IBUF(m1_m1_dataout[20]),.OUT_IBUF(m1_m1_dataout_int[20]));

	qlIBUF QL_INST_A2F_B_20_4 (.IN_IBUF(m1_m1_dataout[19]),.OUT_IBUF(m1_m1_dataout_int[19]));

	qlIBUF QL_INST_A2F_B_20_5 (.IN_IBUF(m1_m1_dataout[18]),.OUT_IBUF(m1_m1_dataout_int[18]));

	qlIBUF QL_INST_A2F_B_20_6 (.IN_IBUF(m1_m1_dataout[17]),.OUT_IBUF(m1_m1_dataout_int[17]));

	qlOBUF QL_INST_F2A_B_21_0 (.IN_OBUF(m1_coef_rdata_int[5]),.OUT_OBUF(m1_m1_coef_in[5]));

	qlOBUF QL_INST_F2A_B_21_1 (.IN_OBUF(m1_coef_rdata_int[4]),.OUT_OBUF(m1_m1_coef_in[4]));

	qlOBUF QL_INST_F2A_B_21_2 (.IN_OBUF(m1_coef_rdata_int[3]),.OUT_OBUF(m1_m1_coef_in[3]));

	qlOBUF QL_INST_F2A_B_21_3 (.IN_OBUF(m1_coef_rdata_int[2]),.OUT_OBUF(m1_m1_coef_in[2]));

	qlOBUF QL_INST_F2A_B_21_4 (.IN_OBUF(m1_coef_rdata_int[1]),.OUT_OBUF(m1_m1_coef_in[1]));

	qlOBUF QL_INST_F2A_B_21_5 (.IN_OBUF(m1_coef_rdata_int[0]),.OUT_OBUF(m1_m1_coef_in[0]));

	qlOBUF QL_INST_F2A_B_21_6 (.IN_OBUF(m1_m1_mode_dup_0[1]),.OUT_OBUF(m1_m1_mode[1]));

	qlOBUF QL_INST_F2A_B_21_7 (.IN_OBUF(m1_m1_csel_dup_0),.OUT_OBUF(m1_m1_csel));

	qlOBUF QL_INST_F2A_B_21_8 (.IN_OBUF(m1_m1_mode_dup_0[0]),.OUT_OBUF(m1_m1_mode[0]));

	qlOBUF QL_INST_F2A_B_21_9 (.IN_OBUF(m1_oper1_rdata_int[31]),.OUT_OBUF(m1_m1_oper_in[31]));

	qlOBUF QL_INST_F2A_B_21_10 (.IN_OBUF(m1_oper1_rdata_int[30]),.OUT_OBUF(m1_m1_oper_in[30]));

	qlOBUF QL_INST_F2A_B_21_11 (.IN_OBUF(m1_oper1_rdata_int[29]),.OUT_OBUF(m1_m1_oper_in[29]));

	qlIBUF QL_INST_A2F_B_21_0 (.IN_IBUF(m1_m1_dataout[16]),.OUT_IBUF(m1_m1_dataout_int[16]));

	qlIBUF QL_INST_A2F_B_21_1 (.IN_IBUF(m1_m1_dataout[15]),.OUT_IBUF(m1_m1_dataout_int[15]));

	qlIBUF QL_INST_A2F_B_21_2 (.IN_IBUF(m1_m1_dataout[14]),.OUT_IBUF(m1_m1_dataout_int[14]));

	qlIBUF QL_INST_A2F_B_21_3 (.IN_IBUF(m1_m1_dataout[13]),.OUT_IBUF(m1_m1_dataout_int[13]));

	qlIBUF QL_INST_A2F_B_21_4 (.IN_IBUF(m1_m1_dataout[12]),.OUT_IBUF(m1_m1_dataout_int[12]));

	qlIBUF QL_INST_A2F_B_21_5 (.IN_IBUF(m1_m1_dataout[11]),.OUT_IBUF(m1_m1_dataout_int[11]));

	qlOBUF QL_INST_F2A_B_22_0 (.IN_OBUF(m1_oper1_rdata_int[28]),.OUT_OBUF(m1_m1_oper_in[28]));

	qlOBUF QL_INST_F2A_B_22_1 (.IN_OBUF(m1_oper1_rdata_int[27]),.OUT_OBUF(m1_m1_oper_in[27]));

	qlOBUF QL_INST_F2A_B_22_2 (.IN_OBUF(m1_oper1_rdata_int[26]),.OUT_OBUF(m1_m1_oper_in[26]));

	qlOBUF QL_INST_F2A_B_22_3 (.IN_OBUF(m1_oper1_rdata_int[25]),.OUT_OBUF(m1_m1_oper_in[25]));

	qlOBUF QL_INST_F2A_B_22_4 (.IN_OBUF(m1_oper1_rdata_int[24]),.OUT_OBUF(m1_m1_oper_in[24]));

	qlOBUF QL_INST_F2A_B_22_5 (.IN_OBUF(m1_oper1_rdata_int[23]),.OUT_OBUF(m1_m1_oper_in[23]));

	qlOBUF QL_INST_F2A_B_22_6 (.IN_OBUF(m1_oper1_rdata_int[22]),.OUT_OBUF(m1_m1_oper_in[22]));

	qlOBUF QL_INST_F2A_B_22_7 (.IN_OBUF(m1_oper1_rdata_int[21]),.OUT_OBUF(m1_m1_oper_in[21]));

	qlOBUF QL_INST_F2A_B_22_8 (.IN_OBUF(m1_oper1_rdata_int[20]),.OUT_OBUF(m1_m1_oper_in[20]));

	qlOBUF QL_INST_F2A_B_22_9 (.IN_OBUF(m1_oper1_rdata_int[19]),.OUT_OBUF(m1_m1_oper_in[19]));

	qlOBUF QL_INST_F2A_B_22_10 (.IN_OBUF(m1_oper1_rdata_int[18]),.OUT_OBUF(m1_m1_oper_in[18]));

	qlOBUF QL_INST_F2A_B_22_11 (.IN_OBUF(m1_oper1_rdata_int[17]),.OUT_OBUF(m1_m1_oper_in[17]));

	qlOBUF QL_INST_F2A_B_22_12 (.IN_OBUF(m1_oper1_rdata_int[16]),.OUT_OBUF(m1_m1_oper_in[16]));

	qlOBUF QL_INST_F2A_B_22_13 (.IN_OBUF(m1_oper1_rdata_int[15]),.OUT_OBUF(m1_m1_oper_in[15]));

	qlOBUF QL_INST_F2A_B_22_14 (.IN_OBUF(m1_oper1_rdata_int[14]),.OUT_OBUF(m1_m1_oper_in[14]));

	qlOBUF QL_INST_F2A_B_22_15 (.IN_OBUF(m1_oper1_rdata_int[13]),.OUT_OBUF(m1_m1_oper_in[13]));

	qlOBUF QL_INST_F2A_B_22_16 (.IN_OBUF(m1_oper1_rdata_int[12]),.OUT_OBUF(m1_m1_oper_in[12]));

	qlOBUF QL_INST_F2A_B_22_17 (.IN_OBUF(m1_oper1_rdata_int[11]),.OUT_OBUF(m1_m1_oper_in[11]));

	qlIBUF QL_INST_A2F_B_22_0 (.IN_IBUF(m1_m1_dataout[10]),.OUT_IBUF(m1_m1_dataout_int[10]));

	qlIBUF QL_INST_A2F_B_22_1 (.IN_IBUF(m1_m1_dataout[9]),.OUT_IBUF(m1_m1_dataout_int[9]));

	qlIBUF QL_INST_A2F_B_22_2 (.IN_IBUF(m1_m1_dataout[8]),.OUT_IBUF(m1_m1_dataout_int[8]));

	qlIBUF QL_INST_A2F_B_22_3 (.IN_IBUF(m1_m1_dataout[7]),.OUT_IBUF(m1_m1_dataout_int[7]));

	qlIBUF QL_INST_A2F_B_22_4 (.IN_IBUF(m1_m1_dataout[6]),.OUT_IBUF(m1_m1_dataout_int[6]));

	qlIBUF QL_INST_A2F_B_22_5 (.IN_IBUF(m1_m1_dataout[5]),.OUT_IBUF(m1_m1_dataout_int[5]));

	qlOBUF QL_INST_F2A_B_23_0 (.IN_OBUF(m1_oper1_rdata_int[10]),.OUT_OBUF(m1_m1_oper_in[10]));

	qlOBUF QL_INST_F2A_B_23_1 (.IN_OBUF(m1_oper1_rdata_int[9]),.OUT_OBUF(m1_m1_oper_in[9]));

	qlOBUF QL_INST_F2A_B_23_2 (.IN_OBUF(m1_oper1_rdata_int[8]),.OUT_OBUF(m1_m1_oper_in[8]));

	qlOBUF QL_INST_F2A_B_23_3 (.IN_OBUF(m1_oper1_rdata_int[7]),.OUT_OBUF(m1_m1_oper_in[7]));

	qlOBUF QL_INST_F2A_B_23_4 (.IN_OBUF(m1_oper1_rdata_int[6]),.OUT_OBUF(m1_m1_oper_in[6]));

	qlOBUF QL_INST_F2A_B_23_5 (.IN_OBUF(m1_oper1_rdata_int[5]),.OUT_OBUF(m1_m1_oper_in[5]));

	qlOBUF QL_INST_F2A_B_23_6 (.IN_OBUF(m1_oper1_rdata_int[4]),.OUT_OBUF(m1_m1_oper_in[4]));

	qlOBUF QL_INST_F2A_B_23_7 (.IN_OBUF(m1_oper1_rdata_int[3]),.OUT_OBUF(m1_m1_oper_in[3]));

	qlOBUF QL_INST_F2A_B_23_8 (.IN_OBUF(m1_oper1_rdata_int[2]),.OUT_OBUF(m1_m1_oper_in[2]));

	qlOBUF QL_INST_F2A_B_23_9 (.IN_OBUF(m1_oper1_rdata_int[1]),.OUT_OBUF(m1_m1_oper_in[1]));

	qlOBUF QL_INST_F2A_B_23_10 (.IN_OBUF(m1_oper1_rdata_int[0]),.OUT_OBUF(m1_m1_oper_in[0]));

	qlIBUF QL_INST_A2F_B_23_0 (.IN_IBUF(m1_m1_dataout[4]),.OUT_IBUF(m1_m1_dataout_int[4]));

	qlIBUF QL_INST_A2F_B_23_1 (.IN_IBUF(m1_m1_dataout[3]),.OUT_IBUF(m1_m1_dataout_int[3]));

	qlIBUF QL_INST_A2F_B_23_2 (.IN_IBUF(m1_m1_dataout[2]),.OUT_IBUF(m1_m1_dataout_int[2]));

	qlIBUF QL_INST_A2F_B_23_3 (.IN_IBUF(m1_m1_dataout[1]),.OUT_IBUF(m1_m1_dataout_int[1]));

	qlIBUF QL_INST_A2F_B_23_4 (.IN_IBUF(m1_m1_dataout[0]),.OUT_IBUF(m1_m1_dataout_int[0]));

	qlOBUF QL_INST_F2A_B_24_16 (.IN_OBUF(m1_oper1_wdata_dup_0[31]),.OUT_OBUF(m1_oper1_wdata[31]));

	qlOBUF QL_INST_F2A_B_24_17 (.IN_OBUF(m1_oper1_wdata_dup_0[30]),.OUT_OBUF(m1_oper1_wdata[30]));

	DBUF QL_INST_F2Adef_B_24_1 (.IN_DBUF(GND),.OUT_DBUF(m0_oper0_powerdn));

	qlOBUF QL_INST_F2A_B_25_0 (.IN_OBUF(m1_oper1_wdata_dup_0[29]),.OUT_OBUF(m1_oper1_wdata[29]));

	qlOBUF QL_INST_F2A_B_25_1 (.IN_OBUF(m1_oper1_wdata_dup_0[28]),.OUT_OBUF(m1_oper1_wdata[28]));

	qlOBUF QL_INST_F2A_B_25_2 (.IN_OBUF(m1_oper1_wdata_dup_0[27]),.OUT_OBUF(m1_oper1_wdata[27]));

	qlOBUF QL_INST_F2A_B_25_3 (.IN_OBUF(m1_oper1_wdata_dup_0[26]),.OUT_OBUF(m1_oper1_wdata[26]));

	qlOBUF QL_INST_F2A_B_25_4 (.IN_OBUF(m1_oper1_wdata_dup_0[25]),.OUT_OBUF(m1_oper1_wdata[25]));

	qlOBUF QL_INST_F2A_B_25_5 (.IN_OBUF(m1_oper1_wdata_dup_0[24]),.OUT_OBUF(m1_oper1_wdata[24]));

	qlOBUF QL_INST_F2A_B_25_6 (.IN_OBUF(m1_oper1_wdata_dup_0[23]),.OUT_OBUF(m1_oper1_wdata[23]));

	qlOBUF QL_INST_F2A_B_25_7 (.IN_OBUF(m1_oper1_wdata_dup_0[22]),.OUT_OBUF(m1_oper1_wdata[22]));

	qlOBUF QL_INST_F2A_B_25_8 (.IN_OBUF(m1_oper1_wdata_dup_0[21]),.OUT_OBUF(m1_oper1_wdata[21]));

	qlOBUF QL_INST_F2A_B_25_9 (.IN_OBUF(m1_oper1_wdata_dup_0[20]),.OUT_OBUF(m1_oper1_wdata[20]));

	qlOBUF QL_INST_F2A_B_25_10 (.IN_OBUF(m1_oper1_wdata_dup_0[19]),.OUT_OBUF(m1_oper1_wdata[19]));

	qlOBUF QL_INST_F2A_B_25_11 (.IN_OBUF(m1_oper1_wdata_dup_0[18]),.OUT_OBUF(m1_oper1_wdata[18]));

	qlIBUF QL_INST_A2F_B_25_1 (.IN_IBUF(m1_oper1_rdata[31]),.OUT_IBUF(m1_oper1_rdata_int[31]));

	qlIBUF QL_INST_A2F_B_25_2 (.IN_IBUF(m1_oper1_rdata[30]),.OUT_IBUF(m1_oper1_rdata_int[30]));

	qlIBUF QL_INST_A2F_B_25_3 (.IN_IBUF(m1_oper1_rdata[29]),.OUT_IBUF(m1_oper1_rdata_int[29]));

	qlIBUF QL_INST_A2F_B_25_4 (.IN_IBUF(m1_oper1_rdata[28]),.OUT_IBUF(m1_oper1_rdata_int[28]));

	qlIBUF QL_INST_A2F_B_25_5 (.IN_IBUF(m1_oper1_rdata[27]),.OUT_IBUF(m1_oper1_rdata_int[27]));

	qlOBUF QL_INST_F2A_B_26_0 (.IN_OBUF(m1_oper1_wdata_dup_0[17]),.OUT_OBUF(m1_oper1_wdata[17]));

	qlOBUF QL_INST_F2A_B_26_1 (.IN_OBUF(m1_oper1_wdata_dup_0[16]),.OUT_OBUF(m1_oper1_wdata[16]));

	qlOBUF QL_INST_F2A_B_26_2 (.IN_OBUF(m1_oper1_wdata_dup_0[15]),.OUT_OBUF(m1_oper1_wdata[15]));

	qlOBUF QL_INST_F2A_B_26_3 (.IN_OBUF(m1_oper1_wdata_dup_0[14]),.OUT_OBUF(m1_oper1_wdata[14]));

	qlOBUF QL_INST_F2A_B_26_4 (.IN_OBUF(m1_oper1_wdata_dup_0[13]),.OUT_OBUF(m1_oper1_wdata[13]));

	qlOBUF QL_INST_F2A_B_26_5 (.IN_OBUF(m1_oper1_wdata_dup_0[12]),.OUT_OBUF(m1_oper1_wdata[12]));

	qlOBUF QL_INST_F2A_B_26_6 (.IN_OBUF(m1_oper1_wdata_dup_0[11]),.OUT_OBUF(m1_oper1_wdata[11]));

	qlOBUF QL_INST_F2A_B_26_7 (.IN_OBUF(m1_oper1_wdata_dup_0[10]),.OUT_OBUF(m1_oper1_wdata[10]));

	qlOBUF QL_INST_F2A_B_26_8 (.IN_OBUF(m1_oper1_wdata_dup_0[9]),.OUT_OBUF(m1_oper1_wdata[9]));

	qlOBUF QL_INST_F2A_B_26_9 (.IN_OBUF(m1_oper1_wdata_dup_0[8]),.OUT_OBUF(m1_oper1_wdata[8]));

	qlOBUF QL_INST_F2A_B_26_10 (.IN_OBUF(m1_oper1_wdata_dup_0[7]),.OUT_OBUF(m1_oper1_wdata[7]));

	qlOBUF QL_INST_F2A_B_26_11 (.IN_OBUF(m1_oper1_wdata_dup_0[6]),.OUT_OBUF(m1_oper1_wdata[6]));

	qlOBUF QL_INST_F2A_B_26_12 (.IN_OBUF(m1_oper1_wdata_dup_0[5]),.OUT_OBUF(m1_oper1_wdata[5]));

	qlOBUF QL_INST_F2A_B_26_13 (.IN_OBUF(m1_oper1_wdata_dup_0[4]),.OUT_OBUF(m1_oper1_wdata[4]));

	qlOBUF QL_INST_F2A_B_26_14 (.IN_OBUF(m1_oper1_wdata_dup_0[3]),.OUT_OBUF(m1_oper1_wdata[3]));

	qlOBUF QL_INST_F2A_B_26_15 (.IN_OBUF(m1_oper1_wdata_dup_0[2]),.OUT_OBUF(m1_oper1_wdata[2]));

	qlOBUF QL_INST_F2A_B_26_16 (.IN_OBUF(m1_oper1_wdata_dup_0[1]),.OUT_OBUF(m1_oper1_wdata[1]));

	qlOBUF QL_INST_F2A_B_26_17 (.IN_OBUF(m1_oper1_wdata_dup_0[0]),.OUT_OBUF(m1_oper1_wdata[0]));

	qlIBUF QL_INST_A2F_B_26_0 (.IN_IBUF(m1_oper1_rdata[26]),.OUT_IBUF(m1_oper1_rdata_int[26]));

	qlIBUF QL_INST_A2F_B_26_1 (.IN_IBUF(m1_oper1_rdata[25]),.OUT_IBUF(m1_oper1_rdata_int[25]));

	qlIBUF QL_INST_A2F_B_26_2 (.IN_IBUF(m1_oper1_rdata[24]),.OUT_IBUF(m1_oper1_rdata_int[24]));

	qlIBUF QL_INST_A2F_B_26_3 (.IN_IBUF(m1_oper1_rdata[23]),.OUT_IBUF(m1_oper1_rdata_int[23]));

	qlIBUF QL_INST_A2F_B_26_4 (.IN_IBUF(m1_oper1_rdata[22]),.OUT_IBUF(m1_oper1_rdata_int[22]));

	qlIBUF QL_INST_A2F_B_26_5 (.IN_IBUF(m1_oper1_rdata[21]),.OUT_IBUF(m1_oper1_rdata_int[21]));

	qlIBUF QL_INST_A2F_B_26_6 (.IN_IBUF(m1_oper1_rdata[20]),.OUT_IBUF(m1_oper1_rdata_int[20]));

	qlIBUF QL_INST_A2F_B_26_7 (.IN_IBUF(m1_oper1_rdata[19]),.OUT_IBUF(m1_oper1_rdata_int[19]));

	qlOBUF QL_INST_F2A_B_27_0 (.IN_OBUF(m1_oper1_waddr_dup_0[11]),.OUT_OBUF(m1_oper1_waddr[11]));

	qlOBUF QL_INST_F2A_B_27_1 (.IN_OBUF(m1_oper1_waddr_dup_0[10]),.OUT_OBUF(m1_oper1_waddr[10]));

	qlOBUF QL_INST_F2A_B_27_2 (.IN_OBUF(m1_oper1_waddr_dup_0[9]),.OUT_OBUF(m1_oper1_waddr[9]));

	qlOBUF QL_INST_F2A_B_27_3 (.IN_OBUF(m1_oper1_waddr_dup_0[8]),.OUT_OBUF(m1_oper1_waddr[8]));

	qlOBUF QL_INST_F2A_B_27_4 (.IN_OBUF(m1_oper1_waddr_dup_0[7]),.OUT_OBUF(m1_oper1_waddr[7]));

	qlOBUF QL_INST_F2A_B_27_5 (.IN_OBUF(m1_oper1_waddr_dup_0[6]),.OUT_OBUF(m1_oper1_waddr[6]));

	qlOBUF QL_INST_F2A_B_27_6 (.IN_OBUF(m1_oper1_waddr_dup_0[5]),.OUT_OBUF(m1_oper1_waddr[5]));

	qlOBUF QL_INST_F2A_B_27_7 (.IN_OBUF(m1_oper1_waddr_dup_0[4]),.OUT_OBUF(m1_oper1_waddr[4]));

	qlOBUF QL_INST_F2A_B_27_8 (.IN_OBUF(m1_oper1_waddr_dup_0[3]),.OUT_OBUF(m1_oper1_waddr[3]));

	qlOBUF QL_INST_F2A_B_27_9 (.IN_OBUF(m1_oper1_waddr_dup_0[2]),.OUT_OBUF(m1_oper1_waddr[2]));

	qlOBUF QL_INST_F2A_B_27_10 (.IN_OBUF(m1_oper1_waddr_dup_0[1]),.OUT_OBUF(m1_oper1_waddr[1]));

	qlOBUF QL_INST_F2A_B_27_11 (.IN_OBUF(m1_oper1_waddr_dup_0[0]),.OUT_OBUF(m1_oper1_waddr[0]));

	qlIBUF QL_INST_A2F_B_27_0 (.IN_IBUF(m1_oper1_rdata[18]),.OUT_IBUF(m1_oper1_rdata_int[18]));

	qlIBUF QL_INST_A2F_B_27_1 (.IN_IBUF(m1_oper1_rdata[17]),.OUT_IBUF(m1_oper1_rdata_int[17]));

	qlIBUF QL_INST_A2F_B_27_2 (.IN_IBUF(m1_oper1_rdata[16]),.OUT_IBUF(m1_oper1_rdata_int[16]));

	qlIBUF QL_INST_A2F_B_27_3 (.IN_IBUF(m1_oper1_rdata[15]),.OUT_IBUF(m1_oper1_rdata_int[15]));

	qlIBUF QL_INST_A2F_B_27_4 (.IN_IBUF(m1_oper1_rdata[14]),.OUT_IBUF(m1_oper1_rdata_int[14]));

	qlIBUF QL_INST_A2F_B_27_5 (.IN_IBUF(m1_oper1_rdata[13]),.OUT_IBUF(m1_oper1_rdata_int[13]));

	qlOBUF QL_INST_F2A_B_28_0 (.IN_OBUF(CLK_int_0__CAND0_BRSBR_28_padClk),.OUT_OBUF(m1_oper1_wclk));

	qlOBUF QL_INST_F2A_B_28_1 (.IN_OBUF(m0_oper1_wmode_dup_0[1]),.OUT_OBUF(m1_oper1_wmode[1]));

	qlOBUF QL_INST_F2A_B_28_2 (.IN_OBUF(m0_oper1_wmode_dup_0[0]),.OUT_OBUF(m1_oper1_wmode[0]));

	qlOBUF QL_INST_F2A_B_28_3 (.IN_OBUF(m0_oper1_wdsel_dup_0),.OUT_OBUF(m1_oper1_wdsel));

	qlOBUF QL_INST_F2A_B_28_4 (.IN_OBUF(m1_oper1_we_dup_0),.OUT_OBUF(m1_oper1_we));

	qlOBUF QL_INST_F2A_B_28_15 (.IN_OBUF(m0_oper1_rmode_dup_0[1]),.OUT_OBUF(m1_oper1_rmode[1]));

	qlOBUF QL_INST_F2A_B_28_16 (.IN_OBUF(m0_oper1_rmode_dup_0[0]),.OUT_OBUF(m1_oper1_rmode[0]));

	qlOBUF QL_INST_F2A_B_28_17 (.IN_OBUF(m1_oper1_raddr_dup_0[11]),.OUT_OBUF(m1_oper1_raddr[11]));

	qlIBUF QL_INST_A2F_B_28_1 (.IN_IBUF(m1_oper1_rdata[12]),.OUT_IBUF(m1_oper1_rdata_int[12]));

	qlIBUF QL_INST_A2F_B_28_2 (.IN_IBUF(m1_oper1_rdata[11]),.OUT_IBUF(m1_oper1_rdata_int[11]));

	qlIBUF QL_INST_A2F_B_28_3 (.IN_IBUF(m1_oper1_rdata[10]),.OUT_IBUF(m1_oper1_rdata_int[10]));

	qlIBUF QL_INST_A2F_B_28_4 (.IN_IBUF(m1_oper1_rdata[9]),.OUT_IBUF(m1_oper1_rdata_int[9]));

	qlIBUF QL_INST_A2F_B_28_5 (.IN_IBUF(m1_oper1_rdata[8]),.OUT_IBUF(m1_oper1_rdata_int[8]));

	qlIBUF QL_INST_A2F_B_28_6 (.IN_IBUF(m1_oper1_rdata[7]),.OUT_IBUF(m1_oper1_rdata_int[7]));

	qlIBUF QL_INST_A2F_B_28_7 (.IN_IBUF(m1_oper1_rdata[6]),.OUT_IBUF(m1_oper1_rdata_int[6]));

	qlOBUF QL_INST_F2A_B_29_0 (.IN_OBUF(CLK_int_0__CAND0_BRSBR_29_padClk),.OUT_OBUF(m1_oper1_rclk));

	qlOBUF QL_INST_F2A_B_29_1 (.IN_OBUF(m1_oper1_raddr_dup_0[10]),.OUT_OBUF(m1_oper1_raddr[10]));

	qlOBUF QL_INST_F2A_B_29_2 (.IN_OBUF(m1_oper1_raddr_dup_0[9]),.OUT_OBUF(m1_oper1_raddr[9]));

	qlOBUF QL_INST_F2A_B_29_3 (.IN_OBUF(m1_oper1_raddr_dup_0[8]),.OUT_OBUF(m1_oper1_raddr[8]));

	qlOBUF QL_INST_F2A_B_29_4 (.IN_OBUF(m1_oper1_raddr_dup_0[7]),.OUT_OBUF(m1_oper1_raddr[7]));

	qlOBUF QL_INST_F2A_B_29_5 (.IN_OBUF(m1_oper1_raddr_dup_0[6]),.OUT_OBUF(m1_oper1_raddr[6]));

	qlOBUF QL_INST_F2A_B_29_6 (.IN_OBUF(m1_oper1_raddr_dup_0[5]),.OUT_OBUF(m1_oper1_raddr[5]));

	qlOBUF QL_INST_F2A_B_29_7 (.IN_OBUF(m1_oper1_raddr_dup_0[4]),.OUT_OBUF(m1_oper1_raddr[4]));

	qlOBUF QL_INST_F2A_B_29_8 (.IN_OBUF(m1_oper1_raddr_dup_0[3]),.OUT_OBUF(m1_oper1_raddr[3]));

	qlOBUF QL_INST_F2A_B_29_9 (.IN_OBUF(m1_oper1_raddr_dup_0[2]),.OUT_OBUF(m1_oper1_raddr[2]));

	qlOBUF QL_INST_F2A_B_29_10 (.IN_OBUF(m1_oper1_raddr_dup_0[1]),.OUT_OBUF(m1_oper1_raddr[1]));

	qlOBUF QL_INST_F2A_B_29_11 (.IN_OBUF(m1_oper1_raddr_dup_0[0]),.OUT_OBUF(m1_oper1_raddr[0]));

	qlIBUF QL_INST_A2F_B_29_0 (.IN_IBUF(m1_oper1_rdata[5]),.OUT_IBUF(m1_oper1_rdata_int[5]));

	qlIBUF QL_INST_A2F_B_29_1 (.IN_IBUF(m1_oper1_rdata[4]),.OUT_IBUF(m1_oper1_rdata_int[4]));

	qlIBUF QL_INST_A2F_B_29_2 (.IN_IBUF(m1_oper1_rdata[3]),.OUT_IBUF(m1_oper1_rdata_int[3]));

	qlIBUF QL_INST_A2F_B_29_3 (.IN_IBUF(m1_oper1_rdata[2]),.OUT_IBUF(m1_oper1_rdata_int[2]));

	qlIBUF QL_INST_A2F_B_29_4 (.IN_IBUF(m1_oper1_rdata[1]),.OUT_IBUF(m1_oper1_rdata_int[1]));

	qlIBUF QL_INST_A2F_B_29_5 (.IN_IBUF(m1_oper1_rdata[0]),.OUT_IBUF(m1_oper1_rdata_int[0]));

	qlOBUF QL_INST_F2A_L_1_0 (.IN_OBUF(fpgaio_out_dup_0[0]),.OUT_OBUF(fpgaio_out[0]));

	qlOBUF QL_INST_F2A_L_1_1 (.IN_OBUF(fpgaio_oe_dup_0[0]),.OUT_OBUF(fpgaio_oe[0]));

	qlOBUF QL_INST_F2A_L_1_2 (.IN_OBUF(fpgaio_out_dup_0[1]),.OUT_OBUF(fpgaio_out[1]));

	qlOBUF QL_INST_F2A_L_1_3 (.IN_OBUF(fpgaio_oe_dup_0[1]),.OUT_OBUF(fpgaio_oe[1]));

	qlOBUF QL_INST_F2A_L_1_4 (.IN_OBUF(fpgaio_out_dup_0[2]),.OUT_OBUF(fpgaio_out[2]));

	qlOBUF QL_INST_F2A_L_1_5 (.IN_OBUF(fpgaio_oe_dup_0[2]),.OUT_OBUF(fpgaio_oe[2]));

	qlOBUF QL_INST_F2A_L_1_6 (.IN_OBUF(fpgaio_out_dup_0[3]),.OUT_OBUF(fpgaio_out[3]));

	qlOBUF QL_INST_F2A_L_1_7 (.IN_OBUF(fpgaio_oe_dup_0[3]),.OUT_OBUF(fpgaio_oe[3]));

	qlOBUF QL_INST_F2A_L_1_8 (.IN_OBUF(fpgaio_in_int[0]),.OUT_OBUF(events_o[0]));

	qlIBUF QL_INST_A2F_L_1_0 (.IN_IBUF(fpgaio_in[0]),.OUT_IBUF(fpgaio_in_int[0]));

	qlIBUF QL_INST_A2F_L_1_1 (.IN_IBUF(fpgaio_in[12]),.OUT_IBUF(fpgaio_in_int[12]));

	qlIBUF QL_INST_A2F_L_1_2 (.IN_IBUF(fpgaio_in[2]),.OUT_IBUF(fpgaio_in_int[2]));

	qlIBUF QL_INST_A2F_L_1_3 (.IN_IBUF(fpgaio_in[3]),.OUT_IBUF(fpgaio_in_int[3]));

	qlOBUF QL_INST_F2A_L_2_0 (.IN_OBUF(fpgaio_out_dup_0[4]),.OUT_OBUF(fpgaio_out[4]));

	qlOBUF QL_INST_F2A_L_2_1 (.IN_OBUF(fpgaio_oe_dup_0[4]),.OUT_OBUF(fpgaio_oe[4]));

	qlOBUF QL_INST_F2A_L_2_2 (.IN_OBUF(fpgaio_out_dup_0[5]),.OUT_OBUF(fpgaio_out[5]));

	qlOBUF QL_INST_F2A_L_2_3 (.IN_OBUF(fpgaio_oe_dup_0[5]),.OUT_OBUF(fpgaio_oe[5]));

	qlOBUF QL_INST_F2A_L_2_4 (.IN_OBUF(fpgaio_out_dup_0[6]),.OUT_OBUF(fpgaio_out[6]));

	qlOBUF QL_INST_F2A_L_2_5 (.IN_OBUF(fpgaio_oe_dup_0[6]),.OUT_OBUF(fpgaio_oe[6]));

	qlOBUF QL_INST_F2A_L_2_6 (.IN_OBUF(fpgaio_out_dup_0[7]),.OUT_OBUF(fpgaio_out[7]));

	qlOBUF QL_INST_F2A_L_2_7 (.IN_OBUF(fpgaio_oe_dup_0[7]),.OUT_OBUF(fpgaio_oe[7]));

	qlOBUF QL_INST_F2A_L_2_8 (.IN_OBUF(fpgaio_in_int[1]),.OUT_OBUF(events_o[1]));

	qlIBUF QL_INST_A2F_L_2_0 (.IN_IBUF(fpgaio_in[4]),.OUT_IBUF(fpgaio_in_int[4]));

	qlIBUF QL_INST_A2F_L_2_1 (.IN_IBUF(fpgaio_in[5]),.OUT_IBUF(fpgaio_in_int[5]));

	qlIBUF QL_INST_A2F_L_2_2 (.IN_IBUF(fpgaio_in[6]),.OUT_IBUF(fpgaio_in_int[6]));

	qlIBUF QL_INST_A2F_L_2_3 (.IN_IBUF(fpgaio_in[7]),.OUT_IBUF(fpgaio_in_int[7]));

	qlOBUF QL_INST_F2A_L_3_0 (.IN_OBUF(fpgaio_out_dup_0[8]),.OUT_OBUF(fpgaio_out[8]));

	qlOBUF QL_INST_F2A_L_3_1 (.IN_OBUF(fpgaio_oe_dup_0[8]),.OUT_OBUF(fpgaio_oe[8]));

	qlOBUF QL_INST_F2A_L_3_2 (.IN_OBUF(fpgaio_out_dup_0[9]),.OUT_OBUF(fpgaio_out[9]));

	qlOBUF QL_INST_F2A_L_3_3 (.IN_OBUF(fpgaio_oe_dup_0[9]),.OUT_OBUF(fpgaio_oe[9]));

	qlOBUF QL_INST_F2A_L_3_4 (.IN_OBUF(fpgaio_out_dup_0[10]),.OUT_OBUF(fpgaio_out[10]));

	qlOBUF QL_INST_F2A_L_3_5 (.IN_OBUF(fpgaio_oe_dup_0[10]),.OUT_OBUF(fpgaio_oe[10]));

	qlOBUF QL_INST_F2A_L_3_6 (.IN_OBUF(fpgaio_out_dup_0[11]),.OUT_OBUF(fpgaio_out[11]));

	qlOBUF QL_INST_F2A_L_3_7 (.IN_OBUF(fpgaio_oe_dup_0[11]),.OUT_OBUF(fpgaio_oe[11]));

	qlOBUF QL_INST_F2A_L_3_8 (.IN_OBUF(fpgaio_in_int[2]),.OUT_OBUF(events_o[2]));

	qlIBUF QL_INST_A2F_L_3_0 (.IN_IBUF(fpgaio_in[8]),.OUT_IBUF(fpgaio_in_int[8]));

	qlIBUF QL_INST_A2F_L_3_1 (.IN_IBUF(fpgaio_in[9]),.OUT_IBUF(fpgaio_in_int[9]));

	qlIBUF QL_INST_A2F_L_3_2 (.IN_IBUF(fpgaio_in[10]),.OUT_IBUF(fpgaio_in_int[10]));

	qlIBUF QL_INST_A2F_L_3_3 (.IN_IBUF(fpgaio_in[11]),.OUT_IBUF(fpgaio_in_int[11]));

	qlOBUF QL_INST_F2A_L_4_0 (.IN_OBUF(fpgaio_out_dup_0[12]),.OUT_OBUF(fpgaio_out[12]));

	qlOBUF QL_INST_F2A_L_4_1 (.IN_OBUF(fpgaio_oe_dup_0[12]),.OUT_OBUF(fpgaio_oe[12]));

	qlOBUF QL_INST_F2A_L_4_2 (.IN_OBUF(fpgaio_out_dup_0[13]),.OUT_OBUF(fpgaio_out[13]));

	qlOBUF QL_INST_F2A_L_4_3 (.IN_OBUF(fpgaio_oe_dup_0[13]),.OUT_OBUF(fpgaio_oe[13]));

	qlOBUF QL_INST_F2A_L_4_4 (.IN_OBUF(fpgaio_out_dup_0[14]),.OUT_OBUF(fpgaio_out[14]));

	qlOBUF QL_INST_F2A_L_4_5 (.IN_OBUF(fpgaio_oe_dup_0[14]),.OUT_OBUF(fpgaio_oe[14]));

	qlOBUF QL_INST_F2A_L_4_6 (.IN_OBUF(fpgaio_out_dup_0[15]),.OUT_OBUF(fpgaio_out[15]));

	qlOBUF QL_INST_F2A_L_4_7 (.IN_OBUF(fpgaio_oe_dup_0[15]),.OUT_OBUF(fpgaio_oe[15]));

	qlOBUF QL_INST_F2A_L_4_8 (.IN_OBUF(fpgaio_in_int[3]),.OUT_OBUF(events_o[3]));

	qlIBUF QL_INST_A2F_L_4_0 (.IN_IBUF(fpgaio_in[13]),.OUT_IBUF(fpgaio_in_int[13]));

	qlIBUF QL_INST_A2F_L_4_1 (.IN_IBUF(fpgaio_in[14]),.OUT_IBUF(fpgaio_in_int[14]));

	qlIBUF QL_INST_A2F_L_4_2 (.IN_IBUF(fpgaio_in[15]),.OUT_IBUF(fpgaio_in_int[15]));

	qlIBUF QL_INST_A2F_L_4_3 (.IN_IBUF(fpgaio_in[16]),.OUT_IBUF(fpgaio_in_int[16]));

	qlOBUF QL_INST_F2A_L_5_0 (.IN_OBUF(fpgaio_out_dup_0[16]),.OUT_OBUF(fpgaio_out[16]));

	qlOBUF QL_INST_F2A_L_5_1 (.IN_OBUF(fpgaio_oe_dup_0[16]),.OUT_OBUF(fpgaio_oe[16]));

	qlOBUF QL_INST_F2A_L_5_2 (.IN_OBUF(fpgaio_out_dup_0[17]),.OUT_OBUF(fpgaio_out[17]));

	qlOBUF QL_INST_F2A_L_5_3 (.IN_OBUF(fpgaio_oe_dup_0[17]),.OUT_OBUF(fpgaio_oe[17]));

	qlOBUF QL_INST_F2A_L_5_4 (.IN_OBUF(fpgaio_out_dup_0[18]),.OUT_OBUF(fpgaio_out[18]));

	qlOBUF QL_INST_F2A_L_5_5 (.IN_OBUF(fpgaio_oe_dup_0[18]),.OUT_OBUF(fpgaio_oe[18]));

	qlOBUF QL_INST_F2A_L_5_6 (.IN_OBUF(fpgaio_out_dup_0[19]),.OUT_OBUF(fpgaio_out[19]));

	qlOBUF QL_INST_F2A_L_5_7 (.IN_OBUF(fpgaio_oe_dup_0[19]),.OUT_OBUF(fpgaio_oe[19]));

	qlOBUF QL_INST_F2A_L_5_8 (.IN_OBUF(fpgaio_in_int[4]),.OUT_OBUF(events_o[4]));

	qlIBUF QL_INST_A2F_L_5_0 (.IN_IBUF(RESET[2]),.OUT_IBUF(RESET_int[2]));

	qlIBUF QL_INST_A2F_L_5_1 (.IN_IBUF(fpgaio_in[17]),.OUT_IBUF(fpgaio_in_int[17]));

	qlIBUF QL_INST_A2F_L_5_2 (.IN_IBUF(fpgaio_in[18]),.OUT_IBUF(fpgaio_in_int[18]));

	qlIBUF QL_INST_A2F_L_5_3 (.IN_IBUF(fpgaio_in[19]),.OUT_IBUF(fpgaio_in_int[19]));

	qlIBUF QL_INST_A2F_L_5_4 (.IN_IBUF(fpgaio_in[1]),.OUT_IBUF(fpgaio_in_int[1]));

	qlOBUF QL_INST_F2A_L_6_0 (.IN_OBUF(fpgaio_out_dup_0[20]),.OUT_OBUF(fpgaio_out[20]));

	qlOBUF QL_INST_F2A_L_6_1 (.IN_OBUF(fpgaio_oe_dup_0[20]),.OUT_OBUF(fpgaio_oe[20]));

	qlOBUF QL_INST_F2A_L_6_2 (.IN_OBUF(fpgaio_out_dup_0[21]),.OUT_OBUF(fpgaio_out[21]));

	qlOBUF QL_INST_F2A_L_6_3 (.IN_OBUF(fpgaio_oe_dup_0[21]),.OUT_OBUF(fpgaio_oe[21]));

	qlOBUF QL_INST_F2A_L_6_4 (.IN_OBUF(fpgaio_out_dup_0[22]),.OUT_OBUF(fpgaio_out[22]));

	qlOBUF QL_INST_F2A_L_6_5 (.IN_OBUF(fpgaio_oe_dup_0[22]),.OUT_OBUF(fpgaio_oe[22]));

	qlOBUF QL_INST_F2A_L_6_6 (.IN_OBUF(fpgaio_out_dup_0[23]),.OUT_OBUF(fpgaio_out[23]));

	qlOBUF QL_INST_F2A_L_6_7 (.IN_OBUF(fpgaio_oe_dup_0[23]),.OUT_OBUF(fpgaio_oe[23]));

	qlOBUF QL_INST_F2A_L_6_8 (.IN_OBUF(fpgaio_in_int[5]),.OUT_OBUF(events_o[5]));

	qlIBUF QL_INST_A2F_L_6_0 (.IN_IBUF(fpgaio_in[20]),.OUT_IBUF(fpgaio_in_int[20]));

	qlIBUF QL_INST_A2F_L_6_1 (.IN_IBUF(fpgaio_in[21]),.OUT_IBUF(fpgaio_in_int[21]));

	qlIBUF QL_INST_A2F_L_6_2 (.IN_IBUF(fpgaio_in[22]),.OUT_IBUF(fpgaio_in_int[22]));

	qlIBUF QL_INST_A2F_L_6_3 (.IN_IBUF(fpgaio_in[23]),.OUT_IBUF(fpgaio_in_int[23]));

	qlOBUF QL_INST_F2A_L_7_0 (.IN_OBUF(fpgaio_out_dup_0[24]),.OUT_OBUF(fpgaio_out[24]));

	qlOBUF QL_INST_F2A_L_7_1 (.IN_OBUF(fpgaio_oe_dup_0[24]),.OUT_OBUF(fpgaio_oe[24]));

	qlOBUF QL_INST_F2A_L_7_2 (.IN_OBUF(fpgaio_out_dup_0[25]),.OUT_OBUF(fpgaio_out[25]));

	qlOBUF QL_INST_F2A_L_7_3 (.IN_OBUF(fpgaio_oe_dup_0[25]),.OUT_OBUF(fpgaio_oe[25]));

	qlOBUF QL_INST_F2A_L_7_4 (.IN_OBUF(fpgaio_out_dup_0[26]),.OUT_OBUF(fpgaio_out[26]));

	qlOBUF QL_INST_F2A_L_7_5 (.IN_OBUF(fpgaio_oe_dup_0[26]),.OUT_OBUF(fpgaio_oe[26]));

	qlOBUF QL_INST_F2A_L_7_6 (.IN_OBUF(fpgaio_out_dup_0[27]),.OUT_OBUF(fpgaio_out[27]));

	qlOBUF QL_INST_F2A_L_7_7 (.IN_OBUF(fpgaio_oe_dup_0[27]),.OUT_OBUF(fpgaio_oe[27]));

	qlOBUF QL_INST_F2A_L_7_8 (.IN_OBUF(fpgaio_in_int[6]),.OUT_OBUF(events_o[6]));

	qlIBUF QL_INST_A2F_L_7_0 (.IN_IBUF(fpgaio_in[24]),.OUT_IBUF(fpgaio_in_int[24]));

	qlIBUF QL_INST_A2F_L_7_1 (.IN_IBUF(fpgaio_in[25]),.OUT_IBUF(fpgaio_in_int[25]));

	qlIBUF QL_INST_A2F_L_7_2 (.IN_IBUF(fpgaio_in[26]),.OUT_IBUF(fpgaio_in_int[26]));

	qlIBUF QL_INST_A2F_L_7_3 (.IN_IBUF(fpgaio_in[27]),.OUT_IBUF(fpgaio_in_int[27]));

	qlOBUF QL_INST_F2A_L_8_0 (.IN_OBUF(fpgaio_out_dup_0[28]),.OUT_OBUF(fpgaio_out[28]));

	qlOBUF QL_INST_F2A_L_8_1 (.IN_OBUF(fpgaio_oe_dup_0[28]),.OUT_OBUF(fpgaio_oe[28]));

	qlOBUF QL_INST_F2A_L_8_2 (.IN_OBUF(fpgaio_out_dup_0[29]),.OUT_OBUF(fpgaio_out[29]));

	qlOBUF QL_INST_F2A_L_8_3 (.IN_OBUF(fpgaio_oe_dup_0[29]),.OUT_OBUF(fpgaio_oe[29]));

	qlOBUF QL_INST_F2A_L_8_4 (.IN_OBUF(fpgaio_out_dup_0[30]),.OUT_OBUF(fpgaio_out[30]));

	qlOBUF QL_INST_F2A_L_8_5 (.IN_OBUF(fpgaio_oe_dup_0[30]),.OUT_OBUF(fpgaio_oe[30]));

	qlOBUF QL_INST_F2A_L_8_6 (.IN_OBUF(fpgaio_out_dup_0[31]),.OUT_OBUF(fpgaio_out[31]));

	qlOBUF QL_INST_F2A_L_8_7 (.IN_OBUF(fpgaio_oe_dup_0[31]),.OUT_OBUF(fpgaio_oe[31]));

	qlOBUF QL_INST_F2A_L_8_8 (.IN_OBUF(fpgaio_in_int[7]),.OUT_OBUF(events_o[7]));

	qlIBUF QL_INST_A2F_L_8_0 (.IN_IBUF(fpgaio_in[28]),.OUT_IBUF(fpgaio_in_int[28]));

	qlIBUF QL_INST_A2F_L_8_1 (.IN_IBUF(fpgaio_in[29]),.OUT_IBUF(fpgaio_in_int[29]));

	qlIBUF QL_INST_A2F_L_8_2 (.IN_IBUF(fpgaio_in[30]),.OUT_IBUF(fpgaio_in_int[30]));

	qlIBUF QL_INST_A2F_L_8_3 (.IN_IBUF(fpgaio_in[31]),.OUT_IBUF(fpgaio_in_int[31]));

	qlOBUF QL_INST_F2A_L_9_0 (.IN_OBUF(fpgaio_out_dup_0[64]),.OUT_OBUF(fpgaio_out[64]));

	qlOBUF QL_INST_F2A_L_9_1 (.IN_OBUF(fpgaio_oe_dup_0[64]),.OUT_OBUF(fpgaio_oe[64]));

	qlOBUF QL_INST_F2A_L_9_2 (.IN_OBUF(fpgaio_out_dup_0[65]),.OUT_OBUF(fpgaio_out[65]));

	qlOBUF QL_INST_F2A_L_9_3 (.IN_OBUF(fpgaio_oe_dup_0[65]),.OUT_OBUF(fpgaio_oe[65]));

	qlOBUF QL_INST_F2A_L_9_4 (.IN_OBUF(fpgaio_out_dup_0[66]),.OUT_OBUF(fpgaio_out[66]));

	qlOBUF QL_INST_F2A_L_9_5 (.IN_OBUF(fpgaio_oe_dup_0[66]),.OUT_OBUF(fpgaio_oe[66]));

	qlOBUF QL_INST_F2A_L_9_6 (.IN_OBUF(fpgaio_out_dup_0[67]),.OUT_OBUF(fpgaio_out[67]));

	qlOBUF QL_INST_F2A_L_9_7 (.IN_OBUF(fpgaio_oe_dup_0[67]),.OUT_OBUF(fpgaio_oe[67]));

	qlIBUF QL_INST_A2F_L_9_0 (.IN_IBUF(fpgaio_in[64]),.OUT_IBUF(fpgaio_in_int[64]));

	qlIBUF QL_INST_A2F_L_9_1 (.IN_IBUF(fpgaio_in[65]),.OUT_IBUF(fpgaio_in_int[65]));

	qlIBUF QL_INST_A2F_L_9_2 (.IN_IBUF(fpgaio_in[66]),.OUT_IBUF(fpgaio_in_int[66]));

	qlIBUF QL_INST_A2F_L_9_3 (.IN_IBUF(fpgaio_in[67]),.OUT_IBUF(fpgaio_in_int[67]));

	qlOBUF QL_INST_F2A_L_10_0 (.IN_OBUF(fpgaio_out_dup_0[68]),.OUT_OBUF(fpgaio_out[68]));

	qlOBUF QL_INST_F2A_L_10_1 (.IN_OBUF(fpgaio_oe_dup_0[68]),.OUT_OBUF(fpgaio_oe[68]));

	qlOBUF QL_INST_F2A_L_10_2 (.IN_OBUF(fpgaio_out_dup_0[69]),.OUT_OBUF(fpgaio_out[69]));

	qlOBUF QL_INST_F2A_L_10_3 (.IN_OBUF(fpgaio_oe_dup_0[69]),.OUT_OBUF(fpgaio_oe[69]));

	qlOBUF QL_INST_F2A_L_10_4 (.IN_OBUF(fpgaio_out_dup_0[70]),.OUT_OBUF(fpgaio_out[70]));

	qlOBUF QL_INST_F2A_L_10_5 (.IN_OBUF(fpgaio_oe_dup_0[70]),.OUT_OBUF(fpgaio_oe[70]));

	qlOBUF QL_INST_F2A_L_10_6 (.IN_OBUF(fpgaio_out_dup_0[71]),.OUT_OBUF(fpgaio_out[71]));

	qlOBUF QL_INST_F2A_L_10_7 (.IN_OBUF(fpgaio_oe_dup_0[71]),.OUT_OBUF(fpgaio_oe[71]));

	qlIBUF QL_INST_A2F_L_10_0 (.IN_IBUF(fpgaio_in[68]),.OUT_IBUF(fpgaio_in_int[68]));

	qlIBUF QL_INST_A2F_L_10_1 (.IN_IBUF(fpgaio_in[69]),.OUT_IBUF(fpgaio_in_int[69]));

	qlIBUF QL_INST_A2F_L_10_2 (.IN_IBUF(fpgaio_in[70]),.OUT_IBUF(fpgaio_in_int[70]));

	qlIBUF QL_INST_A2F_L_10_3 (.IN_IBUF(fpgaio_in[71]),.OUT_IBUF(fpgaio_in_int[71]));

	qlOBUF QL_INST_F2A_L_11_0 (.IN_OBUF(fpgaio_out_dup_0[72]),.OUT_OBUF(fpgaio_out[72]));

	qlOBUF QL_INST_F2A_L_11_1 (.IN_OBUF(fpgaio_oe_dup_0[72]),.OUT_OBUF(fpgaio_oe[72]));

	qlOBUF QL_INST_F2A_L_11_2 (.IN_OBUF(fpgaio_out_dup_0[73]),.OUT_OBUF(fpgaio_out[73]));

	qlOBUF QL_INST_F2A_L_11_3 (.IN_OBUF(fpgaio_oe_dup_0[73]),.OUT_OBUF(fpgaio_oe[73]));

	qlOBUF QL_INST_F2A_L_11_4 (.IN_OBUF(fpgaio_out_dup_0[74]),.OUT_OBUF(fpgaio_out[74]));

	qlOBUF QL_INST_F2A_L_11_5 (.IN_OBUF(fpgaio_oe_dup_0[74]),.OUT_OBUF(fpgaio_oe[74]));

	qlOBUF QL_INST_F2A_L_11_6 (.IN_OBUF(fpgaio_out_dup_0[75]),.OUT_OBUF(fpgaio_out[75]));

	qlOBUF QL_INST_F2A_L_11_7 (.IN_OBUF(fpgaio_oe_dup_0[75]),.OUT_OBUF(fpgaio_oe[75]));

	qlIBUF QL_INST_A2F_L_11_0 (.IN_IBUF(fpgaio_in[72]),.OUT_IBUF(fpgaio_in_int[72]));

	qlIBUF QL_INST_A2F_L_11_1 (.IN_IBUF(fpgaio_in[73]),.OUT_IBUF(fpgaio_in_int[73]));

	qlIBUF QL_INST_A2F_L_11_2 (.IN_IBUF(fpgaio_in[74]),.OUT_IBUF(fpgaio_in_int[74]));

	qlIBUF QL_INST_A2F_L_11_3 (.IN_IBUF(fpgaio_in[75]),.OUT_IBUF(fpgaio_in_int[75]));

	qlOBUF QL_INST_F2A_L_12_0 (.IN_OBUF(fpgaio_out_dup_0[76]),.OUT_OBUF(fpgaio_out[76]));

	qlOBUF QL_INST_F2A_L_12_1 (.IN_OBUF(fpgaio_oe_dup_0[76]),.OUT_OBUF(fpgaio_oe[76]));

	qlOBUF QL_INST_F2A_L_12_2 (.IN_OBUF(fpgaio_out_dup_0[77]),.OUT_OBUF(fpgaio_out[77]));

	qlOBUF QL_INST_F2A_L_12_3 (.IN_OBUF(fpgaio_oe_dup_0[77]),.OUT_OBUF(fpgaio_oe[77]));

	qlOBUF QL_INST_F2A_L_12_4 (.IN_OBUF(fpgaio_out_dup_0[78]),.OUT_OBUF(fpgaio_out[78]));

	qlOBUF QL_INST_F2A_L_12_5 (.IN_OBUF(fpgaio_oe_dup_0[78]),.OUT_OBUF(fpgaio_oe[78]));

	qlOBUF QL_INST_F2A_L_12_6 (.IN_OBUF(fpgaio_out_dup_0[79]),.OUT_OBUF(fpgaio_out[79]));

	qlOBUF QL_INST_F2A_L_12_7 (.IN_OBUF(fpgaio_oe_dup_0[79]),.OUT_OBUF(fpgaio_oe[79]));

	qlIBUF QL_INST_A2F_L_12_0 (.IN_IBUF(fpgaio_in[76]),.OUT_IBUF(fpgaio_in_int[76]));

	qlIBUF QL_INST_A2F_L_12_1 (.IN_IBUF(fpgaio_in[77]),.OUT_IBUF(fpgaio_in_int[77]));

	qlIBUF QL_INST_A2F_L_12_2 (.IN_IBUF(fpgaio_in[78]),.OUT_IBUF(fpgaio_in_int[78]));

	qlIBUF QL_INST_A2F_L_12_3 (.IN_IBUF(fpgaio_in[79]),.OUT_IBUF(fpgaio_in_int[79]));

	qlOBUF QL_INST_F2A_L_16_0 (.IN_OBUF(lint_RDATA_dup_0[0]),.OUT_OBUF(lint_RDATA[0]));

	qlOBUF QL_INST_F2A_L_16_1 (.IN_OBUF(lint_RDATA_dup_0[1]),.OUT_OBUF(lint_RDATA[1]));

	qlOBUF QL_INST_F2A_L_16_2 (.IN_OBUF(lint_RDATA_dup_0[2]),.OUT_OBUF(lint_RDATA[2]));

	qlOBUF QL_INST_F2A_L_16_3 (.IN_OBUF(lint_RDATA_dup_0[3]),.OUT_OBUF(lint_RDATA[3]));

	qlOBUF QL_INST_F2A_L_16_4 (.IN_OBUF(lint_RDATA_dup_0[4]),.OUT_OBUF(lint_RDATA[4]));

	qlOBUF QL_INST_F2A_L_16_5 (.IN_OBUF(lint_RDATA_dup_0[5]),.OUT_OBUF(lint_RDATA[5]));

	qlOBUF QL_INST_F2A_L_16_6 (.IN_OBUF(lint_RDATA_dup_0[6]),.OUT_OBUF(lint_RDATA[6]));

	qlOBUF QL_INST_F2A_L_16_7 (.IN_OBUF(lint_RDATA_dup_0[7]),.OUT_OBUF(lint_RDATA[7]));

	qlIBUF QL_INST_A2F_L_16_0 (.IN_IBUF(lint_WDATA[0]),.OUT_IBUF(lint_WDATA_int[0]));

	qlIBUF QL_INST_A2F_L_16_1 (.IN_IBUF(lint_WDATA[1]),.OUT_IBUF(lint_WDATA_int[1]));

	qlIBUF QL_INST_A2F_L_16_2 (.IN_IBUF(lint_WDATA[2]),.OUT_IBUF(lint_WDATA_int[2]));

	qlIBUF QL_INST_A2F_L_16_3 (.IN_IBUF(lint_WDATA[3]),.OUT_IBUF(lint_WDATA_int[3]));

	qlIBUF QL_INST_A2F_L_16_4 (.IN_IBUF(lint_WDATA[4]),.OUT_IBUF(lint_WDATA_int[4]));

	qlIBUF QL_INST_A2F_L_16_5 (.IN_IBUF(lint_WDATA[5]),.OUT_IBUF(lint_WDATA_int[5]));

	qlIBUF QL_INST_A2F_L_16_6 (.IN_IBUF(lint_WDATA[6]),.OUT_IBUF(lint_WDATA_int[6]));

	qlIBUF QL_INST_A2F_L_16_7 (.IN_IBUF(lint_WDATA[7]),.OUT_IBUF(lint_WDATA_int[7]));

	qlOBUF QL_INST_F2A_L_17_0 (.IN_OBUF(lint_RDATA_dup_0[8]),.OUT_OBUF(lint_RDATA[8]));

	qlOBUF QL_INST_F2A_L_17_1 (.IN_OBUF(lint_RDATA_dup_0[9]),.OUT_OBUF(lint_RDATA[9]));

	qlOBUF QL_INST_F2A_L_17_2 (.IN_OBUF(lint_RDATA_dup_0[10]),.OUT_OBUF(lint_RDATA[10]));

	qlOBUF QL_INST_F2A_L_17_3 (.IN_OBUF(lint_RDATA_dup_0[11]),.OUT_OBUF(lint_RDATA[11]));

	qlOBUF QL_INST_F2A_L_17_4 (.IN_OBUF(lint_RDATA_dup_0[12]),.OUT_OBUF(lint_RDATA[12]));

	qlOBUF QL_INST_F2A_L_17_5 (.IN_OBUF(lint_RDATA_dup_0[13]),.OUT_OBUF(lint_RDATA[13]));

	qlOBUF QL_INST_F2A_L_17_6 (.IN_OBUF(lint_RDATA_dup_0[14]),.OUT_OBUF(lint_RDATA[14]));

	qlOBUF QL_INST_F2A_L_17_7 (.IN_OBUF(lint_RDATA_dup_0[15]),.OUT_OBUF(lint_RDATA[15]));

	qlIBUF QL_INST_A2F_L_17_0 (.IN_IBUF(lint_ADDR[0]),.OUT_IBUF(lint_ADDR_int[0]));

	qlIBUF QL_INST_A2F_L_17_1 (.IN_IBUF(lint_ADDR[1]),.OUT_IBUF(lint_ADDR_int[1]));

	qlIBUF QL_INST_A2F_L_17_2 (.IN_IBUF(lint_ADDR[2]),.OUT_IBUF(lint_ADDR_int[2]));

	qlIBUF QL_INST_A2F_L_17_3 (.IN_IBUF(lint_ADDR[3]),.OUT_IBUF(lint_ADDR_int[3]));

	qlIBUF QL_INST_A2F_L_17_4 (.IN_IBUF(lint_ADDR[4]),.OUT_IBUF(lint_ADDR_int[4]));

	qlIBUF QL_INST_A2F_L_17_5 (.IN_IBUF(lint_ADDR[5]),.OUT_IBUF(lint_ADDR_int[5]));

	qlOBUF QL_INST_F2A_L_18_0 (.IN_OBUF(CLK_int_0__CAND0_BLSTL_0_padClk),.OUT_OBUF(APB_CLK));

	qlOBUF QL_INST_F2A_L_18_1 (.IN_OBUF(lint_RDATA_dup_0[16]),.OUT_OBUF(lint_RDATA[16]));

	qlOBUF QL_INST_F2A_L_18_2 (.IN_OBUF(lint_RDATA_dup_0[17]),.OUT_OBUF(lint_RDATA[17]));

	qlOBUF QL_INST_F2A_L_18_3 (.IN_OBUF(lint_RDATA_dup_0[18]),.OUT_OBUF(lint_RDATA[18]));

	qlOBUF QL_INST_F2A_L_18_4 (.IN_OBUF(lint_RDATA_dup_0[19]),.OUT_OBUF(lint_RDATA[19]));

	qlOBUF QL_INST_F2A_L_18_5 (.IN_OBUF(lint_RDATA_dup_0[20]),.OUT_OBUF(lint_RDATA[20]));

	qlOBUF QL_INST_F2A_L_18_6 (.IN_OBUF(lint_RDATA_dup_0[21]),.OUT_OBUF(lint_RDATA[21]));

	qlOBUF QL_INST_F2A_L_18_7 (.IN_OBUF(lint_RDATA_dup_0[22]),.OUT_OBUF(lint_RDATA[22]));

	qlOBUF QL_INST_F2A_L_18_8 (.IN_OBUF(lint_RDATA_dup_0[23]),.OUT_OBUF(lint_RDATA[23]));

	qlOBUF QL_INST_F2A_L_18_9 (.IN_OBUF(lint_VALID_dup_0),.OUT_OBUF(lint_VALID));

	qlIBUF QL_INST_A2F_L_18_0 (.IN_IBUF(lint_WDATA[8]),.OUT_IBUF(lint_WDATA_int[8]));

	qlIBUF QL_INST_A2F_L_18_1 (.IN_IBUF(lint_WDATA[9]),.OUT_IBUF(lint_WDATA_int[9]));

	qlIBUF QL_INST_A2F_L_18_2 (.IN_IBUF(lint_WDATA[10]),.OUT_IBUF(lint_WDATA_int[10]));

	qlIBUF QL_INST_A2F_L_18_3 (.IN_IBUF(lint_WDATA[11]),.OUT_IBUF(lint_WDATA_int[11]));

	qlIBUF QL_INST_A2F_L_18_4 (.IN_IBUF(lint_WDATA[12]),.OUT_IBUF(lint_WDATA_int[12]));

	qlIBUF QL_INST_A2F_L_18_5 (.IN_IBUF(lint_WDATA[13]),.OUT_IBUF(lint_WDATA_int[13]));

	qlIBUF QL_INST_A2F_L_18_6 (.IN_IBUF(lint_WDATA[14]),.OUT_IBUF(lint_WDATA_int[14]));

	qlIBUF QL_INST_A2F_L_18_7 (.IN_IBUF(lint_WDATA[15]),.OUT_IBUF(lint_WDATA_int[15]));

	qlOBUF QL_INST_F2A_L_19_1 (.IN_OBUF(lint_RDATA_dup_0[24]),.OUT_OBUF(lint_RDATA[24]));

	qlOBUF QL_INST_F2A_L_19_2 (.IN_OBUF(lint_RDATA_dup_0[25]),.OUT_OBUF(lint_RDATA[25]));

	qlOBUF QL_INST_F2A_L_19_3 (.IN_OBUF(lint_RDATA_dup_0[26]),.OUT_OBUF(lint_RDATA[26]));

	qlOBUF QL_INST_F2A_L_19_4 (.IN_OBUF(lint_RDATA_dup_0[27]),.OUT_OBUF(lint_RDATA[27]));

	qlOBUF QL_INST_F2A_L_19_5 (.IN_OBUF(lint_RDATA_dup_0[28]),.OUT_OBUF(lint_RDATA[28]));

	qlOBUF QL_INST_F2A_L_19_6 (.IN_OBUF(lint_RDATA_dup_0[29]),.OUT_OBUF(lint_RDATA[29]));

	qlOBUF QL_INST_F2A_L_19_7 (.IN_OBUF(lint_RDATA_dup_0[30]),.OUT_OBUF(lint_RDATA[30]));

	qlOBUF QL_INST_F2A_L_19_8 (.IN_OBUF(lint_RDATA_dup_0[31]),.OUT_OBUF(lint_RDATA[31]));

	qlOBUF QL_INST_F2A_L_19_9 (.IN_OBUF(lint_GNT_dup_0),.OUT_OBUF(lint_GNT));

	qlIBUF QL_INST_A2F_L_19_0 (.IN_IBUF(lint_ADDR[6]),.OUT_IBUF(lint_ADDR_int[6]));

	qlIBUF QL_INST_A2F_L_19_1 (.IN_IBUF(lint_ADDR[7]),.OUT_IBUF(lint_ADDR_int[7]));

	qlIBUF QL_INST_A2F_L_19_2 (.IN_IBUF(lint_ADDR[8]),.OUT_IBUF(lint_ADDR_int[8]));

	qlIBUF QL_INST_A2F_L_19_3 (.IN_IBUF(lint_ADDR[9]),.OUT_IBUF(lint_ADDR_int[9]));

	qlIBUF QL_INST_A2F_L_19_4 (.IN_IBUF(lint_ADDR[10]),.OUT_IBUF(lint_ADDR_int[10]));

	qlIBUF QL_INST_A2F_L_19_5 (.IN_IBUF(lint_ADDR[11]),.OUT_IBUF(lint_ADDR_int[11]));

	qlIBUF QL_INST_A2F_L_20_0 (.IN_IBUF(lint_WDATA[16]),.OUT_IBUF(lint_WDATA_int[16]));

	qlIBUF QL_INST_A2F_L_20_1 (.IN_IBUF(lint_WDATA[17]),.OUT_IBUF(lint_WDATA_int[17]));

	qlIBUF QL_INST_A2F_L_20_2 (.IN_IBUF(lint_WDATA[18]),.OUT_IBUF(lint_WDATA_int[18]));

	qlIBUF QL_INST_A2F_L_20_3 (.IN_IBUF(lint_WDATA[19]),.OUT_IBUF(lint_WDATA_int[19]));

	qlIBUF QL_INST_A2F_L_20_4 (.IN_IBUF(lint_WDATA[20]),.OUT_IBUF(lint_WDATA_int[20]));

	qlIBUF QL_INST_A2F_L_20_5 (.IN_IBUF(lint_WDATA[21]),.OUT_IBUF(lint_WDATA_int[21]));

	qlIBUF QL_INST_A2F_L_20_6 (.IN_IBUF(lint_WDATA[22]),.OUT_IBUF(lint_WDATA_int[22]));

	qlIBUF QL_INST_A2F_L_20_7 (.IN_IBUF(lint_WDATA[23]),.OUT_IBUF(lint_WDATA_int[23]));

	qlIBUF QL_INST_A2F_L_21_0 (.IN_IBUF(lint_ADDR[12]),.OUT_IBUF(lint_ADDR_int[12]));

	qlIBUF QL_INST_A2F_L_21_1 (.IN_IBUF(lint_ADDR[13]),.OUT_IBUF(lint_ADDR_int[13]));

	qlIBUF QL_INST_A2F_L_21_2 (.IN_IBUF(lint_ADDR[14]),.OUT_IBUF(lint_ADDR_int[14]));

	qlIBUF QL_INST_A2F_L_21_3 (.IN_IBUF(lint_ADDR[15]),.OUT_IBUF(lint_ADDR_int[15]));

	qlIBUF QL_INST_A2F_L_21_4 (.IN_IBUF(lint_ADDR[16]),.OUT_IBUF(lint_ADDR_int[16]));

	qlIBUF QL_INST_A2F_L_21_5 (.IN_IBUF(lint_ADDR[17]),.OUT_IBUF(lint_ADDR_int[17]));

	qlIBUF QL_INST_A2F_L_22_0 (.IN_IBUF(lint_WDATA[24]),.OUT_IBUF(lint_WDATA_int[24]));

	qlIBUF QL_INST_A2F_L_22_1 (.IN_IBUF(lint_WDATA[25]),.OUT_IBUF(lint_WDATA_int[25]));

	qlIBUF QL_INST_A2F_L_22_2 (.IN_IBUF(lint_WDATA[26]),.OUT_IBUF(lint_WDATA_int[26]));

	qlIBUF QL_INST_A2F_L_22_3 (.IN_IBUF(lint_WDATA[27]),.OUT_IBUF(lint_WDATA_int[27]));

	qlIBUF QL_INST_A2F_L_22_4 (.IN_IBUF(lint_WDATA[28]),.OUT_IBUF(lint_WDATA_int[28]));

	qlIBUF QL_INST_A2F_L_22_5 (.IN_IBUF(lint_WDATA[29]),.OUT_IBUF(lint_WDATA_int[29]));

	qlIBUF QL_INST_A2F_L_22_6 (.IN_IBUF(lint_WDATA[30]),.OUT_IBUF(lint_WDATA_int[30]));

	qlIBUF QL_INST_A2F_L_22_7 (.IN_IBUF(lint_WDATA[31]),.OUT_IBUF(lint_WDATA_int[31]));

	qlIBUF QL_INST_A2F_L_23_0 (.IN_IBUF(lint_ADDR[18]),.OUT_IBUF(lint_ADDR_int[18]));

	qlIBUF QL_INST_A2F_L_23_1 (.IN_IBUF(lint_ADDR[19]),.OUT_IBUF(lint_ADDR_int[19]));

	qlIBUF QL_INST_A2F_L_23_2 (.IN_IBUF(lint_REQ),.OUT_IBUF(lint_REQ_int));

	qlIBUF QL_INST_A2F_L_23_3 (.IN_IBUF(lint_WEN),.OUT_IBUF(lint_WEN_int));

	qlIBUF QL_INST_A2F_L_23_4 (.IN_IBUF(lint_BE[0]),.OUT_IBUF(lint_BE_int[0]));

	qlIBUF QL_INST_A2F_L_23_5 (.IN_IBUF(lint_BE[1]),.OUT_IBUF(lint_BE_int[1]));

	qlIBUF QL_INST_A2F_L_24_0 (.IN_IBUF(lint_BE[2]),.OUT_IBUF(lint_BE_int[2]));

	qlIBUF QL_INST_A2F_L_24_1 (.IN_IBUF(lint_BE[3]),.OUT_IBUF(lint_BE_int[3]));

	qlOBUF QL_INST_F2A_L_25_0 (.IN_OBUF(fpgaio_out_dup_0[32]),.OUT_OBUF(fpgaio_out[32]));

	qlOBUF QL_INST_F2A_L_25_1 (.IN_OBUF(fpgaio_oe_dup_0[32]),.OUT_OBUF(fpgaio_oe[32]));

	qlOBUF QL_INST_F2A_L_25_2 (.IN_OBUF(fpgaio_out_dup_0[33]),.OUT_OBUF(fpgaio_out[33]));

	qlOBUF QL_INST_F2A_L_25_3 (.IN_OBUF(fpgaio_oe_dup_0[33]),.OUT_OBUF(fpgaio_oe[33]));

	qlOBUF QL_INST_F2A_L_25_4 (.IN_OBUF(fpgaio_out_dup_0[34]),.OUT_OBUF(fpgaio_out[34]));

	qlOBUF QL_INST_F2A_L_25_5 (.IN_OBUF(fpgaio_oe_dup_0[34]),.OUT_OBUF(fpgaio_oe[34]));

	qlOBUF QL_INST_F2A_L_25_6 (.IN_OBUF(fpgaio_out_dup_0[35]),.OUT_OBUF(fpgaio_out[35]));

	qlOBUF QL_INST_F2A_L_25_7 (.IN_OBUF(fpgaio_oe_dup_0[35]),.OUT_OBUF(fpgaio_oe[35]));

	qlOBUF QL_INST_F2A_L_25_8 (.IN_OBUF(fpgaio_in_int[8]),.OUT_OBUF(events_o[8]));

	qlIBUF QL_INST_A2F_L_25_0 (.IN_IBUF(fpgaio_in[32]),.OUT_IBUF(fpgaio_in_int[32]));

	qlIBUF QL_INST_A2F_L_25_1 (.IN_IBUF(fpgaio_in[33]),.OUT_IBUF(fpgaio_in_int[33]));

	qlIBUF QL_INST_A2F_L_25_2 (.IN_IBUF(RESET[3]),.OUT_IBUF(RESET_int[3]));

	qlIBUF QL_INST_A2F_L_25_3 (.IN_IBUF(fpgaio_in[34]),.OUT_IBUF(fpgaio_in_int[34]));

	qlIBUF QL_INST_A2F_L_25_4 (.IN_IBUF(fpgaio_in[35]),.OUT_IBUF(fpgaio_in_int[35]));

	qlOBUF QL_INST_F2A_L_26_0 (.IN_OBUF(fpgaio_out_dup_0[36]),.OUT_OBUF(fpgaio_out[36]));

	qlOBUF QL_INST_F2A_L_26_1 (.IN_OBUF(fpgaio_oe_dup_0[36]),.OUT_OBUF(fpgaio_oe[36]));

	qlOBUF QL_INST_F2A_L_26_2 (.IN_OBUF(fpgaio_out_dup_0[37]),.OUT_OBUF(fpgaio_out[37]));

	qlOBUF QL_INST_F2A_L_26_3 (.IN_OBUF(fpgaio_oe_dup_0[37]),.OUT_OBUF(fpgaio_oe[37]));

	qlOBUF QL_INST_F2A_L_26_4 (.IN_OBUF(fpgaio_out_dup_0[38]),.OUT_OBUF(fpgaio_out[38]));

	qlOBUF QL_INST_F2A_L_26_5 (.IN_OBUF(fpgaio_oe_dup_0[38]),.OUT_OBUF(fpgaio_oe[38]));

	qlOBUF QL_INST_F2A_L_26_6 (.IN_OBUF(fpgaio_out_dup_0[39]),.OUT_OBUF(fpgaio_out[39]));

	qlOBUF QL_INST_F2A_L_26_7 (.IN_OBUF(fpgaio_oe_dup_0[39]),.OUT_OBUF(fpgaio_oe[39]));

	qlOBUF QL_INST_F2A_L_26_8 (.IN_OBUF(fpgaio_in_int[9]),.OUT_OBUF(events_o[9]));

	qlIBUF QL_INST_A2F_L_26_0 (.IN_IBUF(fpgaio_in[36]),.OUT_IBUF(fpgaio_in_int[36]));

	qlIBUF QL_INST_A2F_L_26_1 (.IN_IBUF(fpgaio_in[37]),.OUT_IBUF(fpgaio_in_int[37]));

	qlIBUF QL_INST_A2F_L_26_2 (.IN_IBUF(fpgaio_in[38]),.OUT_IBUF(fpgaio_in_int[38]));

	qlIBUF QL_INST_A2F_L_26_3 (.IN_IBUF(fpgaio_in[39]),.OUT_IBUF(fpgaio_in_int[39]));

	qlOBUF QL_INST_F2A_L_27_0 (.IN_OBUF(fpgaio_out_dup_0[40]),.OUT_OBUF(fpgaio_out[40]));

	qlOBUF QL_INST_F2A_L_27_1 (.IN_OBUF(fpgaio_oe_dup_0[40]),.OUT_OBUF(fpgaio_oe[40]));

	qlOBUF QL_INST_F2A_L_27_2 (.IN_OBUF(fpgaio_out_dup_0[41]),.OUT_OBUF(fpgaio_out[41]));

	qlOBUF QL_INST_F2A_L_27_3 (.IN_OBUF(fpgaio_oe_dup_0[41]),.OUT_OBUF(fpgaio_oe[41]));

	qlOBUF QL_INST_F2A_L_27_4 (.IN_OBUF(fpgaio_out_dup_0[42]),.OUT_OBUF(fpgaio_out[42]));

	qlOBUF QL_INST_F2A_L_27_5 (.IN_OBUF(fpgaio_oe_dup_0[42]),.OUT_OBUF(fpgaio_oe[42]));

	qlOBUF QL_INST_F2A_L_27_6 (.IN_OBUF(fpgaio_out_dup_0[43]),.OUT_OBUF(fpgaio_out[43]));

	qlOBUF QL_INST_F2A_L_27_7 (.IN_OBUF(fpgaio_oe_dup_0[43]),.OUT_OBUF(fpgaio_oe[43]));

	qlOBUF QL_INST_F2A_L_27_8 (.IN_OBUF(fpgaio_in_int[10]),.OUT_OBUF(events_o[10]));

	qlIBUF QL_INST_A2F_L_27_0 (.IN_IBUF(fpgaio_in[40]),.OUT_IBUF(fpgaio_in_int[40]));

	qlIBUF QL_INST_A2F_L_27_1 (.IN_IBUF(fpgaio_in[41]),.OUT_IBUF(fpgaio_in_int[41]));

	qlIBUF QL_INST_A2F_L_27_2 (.IN_IBUF(fpgaio_in[42]),.OUT_IBUF(fpgaio_in_int[42]));

	qlIBUF QL_INST_A2F_L_27_3 (.IN_IBUF(fpgaio_in[43]),.OUT_IBUF(fpgaio_in_int[43]));

	qlOBUF QL_INST_F2A_L_28_0 (.IN_OBUF(fpgaio_out_dup_0[44]),.OUT_OBUF(fpgaio_out[44]));

	qlOBUF QL_INST_F2A_L_28_1 (.IN_OBUF(fpgaio_oe_dup_0[44]),.OUT_OBUF(fpgaio_oe[44]));

	qlOBUF QL_INST_F2A_L_28_2 (.IN_OBUF(fpgaio_out_dup_0[45]),.OUT_OBUF(fpgaio_out[45]));

	qlOBUF QL_INST_F2A_L_28_3 (.IN_OBUF(fpgaio_oe_dup_0[45]),.OUT_OBUF(fpgaio_oe[45]));

	qlOBUF QL_INST_F2A_L_28_4 (.IN_OBUF(fpgaio_out_dup_0[46]),.OUT_OBUF(fpgaio_out[46]));

	qlOBUF QL_INST_F2A_L_28_5 (.IN_OBUF(fpgaio_oe_dup_0[46]),.OUT_OBUF(fpgaio_oe[46]));

	qlOBUF QL_INST_F2A_L_28_6 (.IN_OBUF(fpgaio_out_dup_0[47]),.OUT_OBUF(fpgaio_out[47]));

	qlOBUF QL_INST_F2A_L_28_7 (.IN_OBUF(fpgaio_oe_dup_0[47]),.OUT_OBUF(fpgaio_oe[47]));

	qlOBUF QL_INST_F2A_L_28_8 (.IN_OBUF(fpgaio_in_int[11]),.OUT_OBUF(events_o[11]));

	qlIBUF QL_INST_A2F_L_28_0 (.IN_IBUF(fpgaio_in[44]),.OUT_IBUF(fpgaio_in_int[44]));

	qlIBUF QL_INST_A2F_L_28_1 (.IN_IBUF(fpgaio_in[45]),.OUT_IBUF(fpgaio_in_int[45]));

	qlIBUF QL_INST_A2F_L_28_2 (.IN_IBUF(fpgaio_in[46]),.OUT_IBUF(fpgaio_in_int[46]));

	qlIBUF QL_INST_A2F_L_28_3 (.IN_IBUF(fpgaio_in[47]),.OUT_IBUF(fpgaio_in_int[47]));

	qlOBUF QL_INST_F2A_L_29_0 (.IN_OBUF(fpgaio_out_dup_0[48]),.OUT_OBUF(fpgaio_out[48]));

	qlOBUF QL_INST_F2A_L_29_1 (.IN_OBUF(fpgaio_oe_dup_0[48]),.OUT_OBUF(fpgaio_oe[48]));

	qlOBUF QL_INST_F2A_L_29_2 (.IN_OBUF(fpgaio_out_dup_0[49]),.OUT_OBUF(fpgaio_out[49]));

	qlOBUF QL_INST_F2A_L_29_3 (.IN_OBUF(fpgaio_oe_dup_0[49]),.OUT_OBUF(fpgaio_oe[49]));

	qlOBUF QL_INST_F2A_L_29_4 (.IN_OBUF(fpgaio_out_dup_0[50]),.OUT_OBUF(fpgaio_out[50]));

	qlOBUF QL_INST_F2A_L_29_5 (.IN_OBUF(fpgaio_oe_dup_0[50]),.OUT_OBUF(fpgaio_oe[50]));

	qlOBUF QL_INST_F2A_L_29_6 (.IN_OBUF(fpgaio_out_dup_0[51]),.OUT_OBUF(fpgaio_out[51]));

	qlOBUF QL_INST_F2A_L_29_7 (.IN_OBUF(fpgaio_oe_dup_0[51]),.OUT_OBUF(fpgaio_oe[51]));

	qlOBUF QL_INST_F2A_L_29_8 (.IN_OBUF(fpgaio_in_int[12]),.OUT_OBUF(events_o[12]));

	qlIBUF QL_INST_A2F_L_29_0 (.IN_IBUF(fpgaio_in[48]),.OUT_IBUF(fpgaio_in_int[48]));

	qlIBUF QL_INST_A2F_L_29_1 (.IN_IBUF(fpgaio_in[49]),.OUT_IBUF(fpgaio_in_int[49]));

	qlIBUF QL_INST_A2F_L_29_2 (.IN_IBUF(fpgaio_in[50]),.OUT_IBUF(fpgaio_in_int[50]));

	qlIBUF QL_INST_A2F_L_29_3 (.IN_IBUF(fpgaio_in[51]),.OUT_IBUF(fpgaio_in_int[51]));

	qlOBUF QL_INST_F2A_L_30_0 (.IN_OBUF(fpgaio_out_dup_0[52]),.OUT_OBUF(fpgaio_out[52]));

	qlOBUF QL_INST_F2A_L_30_1 (.IN_OBUF(fpgaio_oe_dup_0[52]),.OUT_OBUF(fpgaio_oe[52]));

	qlOBUF QL_INST_F2A_L_30_2 (.IN_OBUF(fpgaio_out_dup_0[53]),.OUT_OBUF(fpgaio_out[53]));

	qlOBUF QL_INST_F2A_L_30_3 (.IN_OBUF(fpgaio_oe_dup_0[53]),.OUT_OBUF(fpgaio_oe[53]));

	qlOBUF QL_INST_F2A_L_30_4 (.IN_OBUF(fpgaio_out_dup_0[54]),.OUT_OBUF(fpgaio_out[54]));

	qlOBUF QL_INST_F2A_L_30_5 (.IN_OBUF(fpgaio_oe_dup_0[54]),.OUT_OBUF(fpgaio_oe[54]));

	qlOBUF QL_INST_F2A_L_30_6 (.IN_OBUF(fpgaio_out_dup_0[55]),.OUT_OBUF(fpgaio_out[55]));

	qlOBUF QL_INST_F2A_L_30_7 (.IN_OBUF(fpgaio_oe_dup_0[55]),.OUT_OBUF(fpgaio_oe[55]));

	qlOBUF QL_INST_F2A_L_30_8 (.IN_OBUF(fpgaio_in_int[13]),.OUT_OBUF(events_o[13]));

	qlIBUF QL_INST_A2F_L_30_0 (.IN_IBUF(fpgaio_in[52]),.OUT_IBUF(fpgaio_in_int[52]));

	qlIBUF QL_INST_A2F_L_30_1 (.IN_IBUF(fpgaio_in[53]),.OUT_IBUF(fpgaio_in_int[53]));

	qlIBUF QL_INST_A2F_L_30_2 (.IN_IBUF(fpgaio_in[54]),.OUT_IBUF(fpgaio_in_int[54]));

	qlIBUF QL_INST_A2F_L_30_3 (.IN_IBUF(fpgaio_in[55]),.OUT_IBUF(fpgaio_in_int[55]));

	qlOBUF QL_INST_F2A_L_31_0 (.IN_OBUF(fpgaio_out_dup_0[56]),.OUT_OBUF(fpgaio_out[56]));

	qlOBUF QL_INST_F2A_L_31_1 (.IN_OBUF(fpgaio_oe_dup_0[56]),.OUT_OBUF(fpgaio_oe[56]));

	qlOBUF QL_INST_F2A_L_31_2 (.IN_OBUF(fpgaio_out_dup_0[57]),.OUT_OBUF(fpgaio_out[57]));

	qlOBUF QL_INST_F2A_L_31_3 (.IN_OBUF(fpgaio_oe_dup_0[57]),.OUT_OBUF(fpgaio_oe[57]));

	qlOBUF QL_INST_F2A_L_31_4 (.IN_OBUF(fpgaio_out_dup_0[58]),.OUT_OBUF(fpgaio_out[58]));

	qlOBUF QL_INST_F2A_L_31_5 (.IN_OBUF(fpgaio_oe_dup_0[58]),.OUT_OBUF(fpgaio_oe[58]));

	qlOBUF QL_INST_F2A_L_31_6 (.IN_OBUF(fpgaio_out_dup_0[59]),.OUT_OBUF(fpgaio_out[59]));

	qlOBUF QL_INST_F2A_L_31_7 (.IN_OBUF(fpgaio_oe_dup_0[59]),.OUT_OBUF(fpgaio_oe[59]));

	qlOBUF QL_INST_F2A_L_31_8 (.IN_OBUF(fpgaio_in_int[14]),.OUT_OBUF(events_o[14]));

	qlIBUF QL_INST_A2F_L_31_0 (.IN_IBUF(fpgaio_in[56]),.OUT_IBUF(fpgaio_in_int[56]));

	qlIBUF QL_INST_A2F_L_31_1 (.IN_IBUF(fpgaio_in[57]),.OUT_IBUF(fpgaio_in_int[57]));

	qlIBUF QL_INST_A2F_L_31_2 (.IN_IBUF(fpgaio_in[58]),.OUT_IBUF(fpgaio_in_int[58]));

	qlIBUF QL_INST_A2F_L_31_3 (.IN_IBUF(fpgaio_in[59]),.OUT_IBUF(fpgaio_in_int[59]));

	qlOBUF QL_INST_F2A_L_32_0 (.IN_OBUF(fpgaio_out_dup_0[60]),.OUT_OBUF(fpgaio_out[60]));

	qlOBUF QL_INST_F2A_L_32_1 (.IN_OBUF(fpgaio_oe_dup_0[60]),.OUT_OBUF(fpgaio_oe[60]));

	qlOBUF QL_INST_F2A_L_32_2 (.IN_OBUF(fpgaio_out_dup_0[61]),.OUT_OBUF(fpgaio_out[61]));

	qlOBUF QL_INST_F2A_L_32_3 (.IN_OBUF(fpgaio_oe_dup_0[61]),.OUT_OBUF(fpgaio_oe[61]));

	qlOBUF QL_INST_F2A_L_32_4 (.IN_OBUF(fpgaio_out_dup_0[62]),.OUT_OBUF(fpgaio_out[62]));

	qlOBUF QL_INST_F2A_L_32_5 (.IN_OBUF(fpgaio_oe_dup_0[62]),.OUT_OBUF(fpgaio_oe[62]));

	qlOBUF QL_INST_F2A_L_32_6 (.IN_OBUF(fpgaio_out_dup_0[63]),.OUT_OBUF(fpgaio_out[63]));

	qlOBUF QL_INST_F2A_L_32_7 (.IN_OBUF(fpgaio_oe_dup_0[63]),.OUT_OBUF(fpgaio_oe[63]));

	qlOBUF QL_INST_F2A_L_32_8 (.IN_OBUF(fpgaio_in_int[15]),.OUT_OBUF(events_o[15]));

	qlIBUF QL_INST_A2F_L_32_0 (.IN_IBUF(fpgaio_in[60]),.OUT_IBUF(fpgaio_in_int[60]));

	qlIBUF QL_INST_A2F_L_32_1 (.IN_IBUF(fpgaio_in[61]),.OUT_IBUF(fpgaio_in_int[61]));

	qlIBUF QL_INST_A2F_L_32_2 (.IN_IBUF(fpgaio_in[62]),.OUT_IBUF(fpgaio_in_int[62]));

	qlIBUF QL_INST_A2F_L_32_3 (.IN_IBUF(fpgaio_in[63]),.OUT_IBUF(fpgaio_in_int[63]));

endmodule


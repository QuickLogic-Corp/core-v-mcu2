/*****************************************************************
          Vendor       : QuickLogic Corp.
          File Name    : top.vq
          Author       : QuickLogic Corp.

          Description : Verilog Simulation Netlist file
******************************************************************/

`timescale 1ns / 10ps

module top1( CLK, RESET, control_in, events_o, fpgaio_in, fpgaio_oe, fpgaio_out, lint_ADDR, lint_BE, lint_GNT, lint_RDATA, lint_REQ, lint_VALID, lint_WDATA, lint_WEN, lint_clk, m0_coef_powerdn, m0_coef_raddr, m0_coef_rclk, m0_coef_rdata, m0_coef_rmode, m0_coef_waddr, m0_coef_wclk, m0_coef_wdata, m0_coef_wdsel, m0_coef_we, m0_coef_wmode, m0_m0_clk, m0_m0_clken, m0_m0_clr, m0_m0_coef_in, m0_m0_csel, m0_m0_dataout, m0_m0_mode, m0_m0_oper_in, m0_m0_osel, m0_m0_outsel, m0_m0_reset, m0_m0_rnd, m0_m0_sat, m0_m0_tc, m0_m1_clk, m0_m1_clken, m0_m1_clr, m0_m1_coef_in, m0_m1_csel, m0_m1_dataout, m0_m1_mode, m0_m1_oper_in, m0_m1_osel, m0_m1_outsel, m0_m1_reset, m0_m1_rnd, m0_m1_sat, m0_m1_tc, m0_oper0_powerdn, m0_oper0_raddr, m0_oper0_rclk, m0_oper0_rdata, m0_oper0_rmode, m0_oper0_waddr, m0_oper0_wclk, m0_oper0_wdata, m0_oper0_wdsel, m0_oper0_we, m0_oper0_wmode, m0_oper1_powerdn, m0_oper1_raddr, m0_oper1_rclk, m0_oper1_rdata, m0_oper1_rmode, m0_oper1_waddr, m0_oper1_wclk, m0_oper1_wdata, m0_oper1_wdsel, m0_oper1_we, m0_oper1_wmode, m1_coef_powerdn, m1_coef_raddr, m1_coef_rclk, m1_coef_rdata, m1_coef_rmode, m1_coef_waddr, m1_coef_wclk, m1_coef_wdata, m1_coef_wdsel, m1_coef_we, m1_coef_wmode, m1_m0_clk, m1_m0_clken, m1_m0_clr, m1_m0_coef_in, m1_m0_csel, m1_m0_dataout, m1_m0_mode, m1_m0_oper_in, m1_m0_osel, m1_m0_outsel, m1_m0_reset, m1_m0_rnd, m1_m0_sat, m1_m0_tc, m1_m1_clk, m1_m1_clken, m1_m1_clr, m1_m1_coef_in, m1_m1_csel, m1_m1_dataout, m1_m1_mode, m1_m1_oper_in, m1_m1_osel, m1_m1_outsel, m1_m1_reset, m1_m1_rnd, m1_m1_sat, m1_m1_tc, m1_oper0_powerdn, m1_oper0_raddr, m1_oper0_rclk, m1_oper0_rdata, m1_oper0_rmode, m1_oper0_waddr, m1_oper0_wclk, m1_oper0_wdata, m1_oper0_wdsel, m1_oper0_we, m1_oper0_wmode, m1_oper1_powerdn, m1_oper1_raddr, m1_oper1_rclk, m1_oper1_rdata, m1_oper1_rmode, m1_oper1_waddr, m1_oper1_wclk, m1_oper1_wdata, m1_oper1_wdsel, m1_oper1_we, m1_oper1_wmode, status_out, tcdm_addr_p0, tcdm_addr_p1, tcdm_addr_p2, tcdm_addr_p3, tcdm_be_p0, tcdm_be_p1, tcdm_be_p2, tcdm_be_p3, tcdm_clk_p0, tcdm_clk_p1, tcdm_clk_p2, tcdm_clk_p3, tcdm_fmo_p0, tcdm_fmo_p1, tcdm_fmo_p2, tcdm_fmo_p3, tcdm_gnt_p0, tcdm_gnt_p1, tcdm_gnt_p2, tcdm_gnt_p3, tcdm_rdata_p0, tcdm_rdata_p1, tcdm_rdata_p2, tcdm_rdata_p3, tcdm_req_p0, tcdm_req_p1, tcdm_req_p2, tcdm_req_p3, tcdm_valid_p0, tcdm_valid_p1, tcdm_valid_p2, tcdm_valid_p3, tcdm_wdata_p0, tcdm_wdata_p1, tcdm_wdata_p2, tcdm_wdata_p3, tcdm_wen_p0, tcdm_wen_p1, tcdm_wen_p2, tcdm_wen_p3, version);
input [5:0] CLK;
input [3:0] RESET;
input [31:0] control_in;
output [15:0] events_o;
input [79:0] fpgaio_in;
output [79:0] fpgaio_oe;
output [79:0] fpgaio_out;
input [19:0] lint_ADDR;
input [3:0] lint_BE;
output lint_GNT;
output [31:0] lint_RDATA;
input lint_REQ;
output lint_VALID;
input [31:0] lint_WDATA;
input lint_WEN;
output lint_clk;
output m0_coef_powerdn;
output [11:0] m0_coef_raddr;
output m0_coef_rclk;
input [31:0] m0_coef_rdata;
output [1:0] m0_coef_rmode;
output [11:0] m0_coef_waddr;
output m0_coef_wclk;
output [31:0] m0_coef_wdata;
output m0_coef_wdsel;
output m0_coef_we;
output [1:0] m0_coef_wmode;
output m0_m0_clk;
output m0_m0_clken;
output m0_m0_clr;
output [31:0] m0_m0_coef_in;
output m0_m0_csel;
input [31:0] m0_m0_dataout;
output [1:0] m0_m0_mode;
output [31:0] m0_m0_oper_in;
output m0_m0_osel;
output [5:0] m0_m0_outsel;
output m0_m0_reset;
output m0_m0_rnd;
output m0_m0_sat;
output m0_m0_tc;
output m0_m1_clk;
output m0_m1_clken;
output m0_m1_clr;
output [31:0] m0_m1_coef_in;
output m0_m1_csel;
input [31:0] m0_m1_dataout;
output [1:0] m0_m1_mode;
output [31:0] m0_m1_oper_in;
output m0_m1_osel;
output [5:0] m0_m1_outsel;
output m0_m1_reset;
output m0_m1_rnd;
output m0_m1_sat;
output m0_m1_tc;
output m0_oper0_powerdn;
output [11:0] m0_oper0_raddr;
output m0_oper0_rclk;
input [31:0] m0_oper0_rdata;
output [1:0] m0_oper0_rmode;
output [11:0] m0_oper0_waddr;
output m0_oper0_wclk;
output [31:0] m0_oper0_wdata;
output m0_oper0_wdsel;
output m0_oper0_we;
output [1:0] m0_oper0_wmode;
output m0_oper1_powerdn;
output [11:0] m0_oper1_raddr;
output m0_oper1_rclk;
input [31:0] m0_oper1_rdata;
output [1:0] m0_oper1_rmode;
output [11:0] m0_oper1_waddr;
output m0_oper1_wclk;
output [31:0] m0_oper1_wdata;
output m0_oper1_wdsel;
output m0_oper1_we;
output [1:0] m0_oper1_wmode;
output m1_coef_powerdn;
output [11:0] m1_coef_raddr;
output m1_coef_rclk;
input [31:0] m1_coef_rdata;
output [1:0] m1_coef_rmode;
output [11:0] m1_coef_waddr;
output m1_coef_wclk;
output [31:0] m1_coef_wdata;
output m1_coef_wdsel;
output m1_coef_we;
output [1:0] m1_coef_wmode;
output m1_m0_clk;
output m1_m0_clken;
output m1_m0_clr;
output [31:0] m1_m0_coef_in;
output m1_m0_csel;
input [31:0] m1_m0_dataout;
output [1:0] m1_m0_mode;
output [31:0] m1_m0_oper_in;
output m1_m0_osel;
output [5:0] m1_m0_outsel;
output m1_m0_reset;
output m1_m0_rnd;
output m1_m0_sat;
output m1_m0_tc;
output m1_m1_clk;
output m1_m1_clken;
output m1_m1_clr;
output [31:0] m1_m1_coef_in;
output m1_m1_csel;
input [31:0] m1_m1_dataout;
output [1:0] m1_m1_mode;
output [31:0] m1_m1_oper_in;
output m1_m1_osel;
output [5:0] m1_m1_outsel;
output m1_m1_reset;
output m1_m1_rnd;
output m1_m1_sat;
output m1_m1_tc;
output m1_oper0_powerdn;
output [11:0] m1_oper0_raddr;
output m1_oper0_rclk;
input [31:0] m1_oper0_rdata;
output [1:0] m1_oper0_rmode;
output [11:0] m1_oper0_waddr;
output m1_oper0_wclk;
output [31:0] m1_oper0_wdata;
output m1_oper0_wdsel;
output m1_oper0_we;
output [1:0] m1_oper0_wmode;
output m1_oper1_powerdn;
output [11:0] m1_oper1_raddr;
output m1_oper1_rclk;
input [31:0] m1_oper1_rdata;
output [1:0] m1_oper1_rmode;
output [11:0] m1_oper1_waddr;
output m1_oper1_wclk;
output [31:0] m1_oper1_wdata;
output m1_oper1_wdsel;
output m1_oper1_we;
output [1:0] m1_oper1_wmode;
output [31:0] status_out;
output [19:0] tcdm_addr_p0;
output [19:0] tcdm_addr_p1;
output [19:0] tcdm_addr_p2;
output [19:0] tcdm_addr_p3;
output [3:0] tcdm_be_p0;
output [3:0] tcdm_be_p1;
output [3:0] tcdm_be_p2;
output [3:0] tcdm_be_p3;
output tcdm_clk_p0;
output tcdm_clk_p1;
output tcdm_clk_p2;
output tcdm_clk_p3;
input tcdm_fmo_p0;
input tcdm_fmo_p1;
input tcdm_fmo_p2;
input tcdm_fmo_p3;
input tcdm_gnt_p0;
input tcdm_gnt_p1;
input tcdm_gnt_p2;
input tcdm_gnt_p3;
input [31:0] tcdm_rdata_p0;
input [31:0] tcdm_rdata_p1;
input [31:0] tcdm_rdata_p2;
input [31:0] tcdm_rdata_p3;
output tcdm_req_p0;
output tcdm_req_p1;
output tcdm_req_p2;
output tcdm_req_p3;
input tcdm_valid_p0;
input tcdm_valid_p1;
input tcdm_valid_p2;
input tcdm_valid_p3;
output [31:0] tcdm_wdata_p0;
output [31:0] tcdm_wdata_p1;
output [31:0] tcdm_wdata_p2;
output [31:0] tcdm_wdata_p3;
output tcdm_wen_p0;
output tcdm_wen_p1;
output tcdm_wen_p2;
output tcdm_wen_p3;
output [7:0] version;

supply1 VCC;
supply0 GND;

wire CLK_int_0__CAND0_BLSBL_1_padClk;
wire CLK_int_0__CAND0_BLSBL_2_padClk;
wire CLK_int_0__CAND0_BLSBL_5_padClk;
wire CLK_int_0__CAND0_BLSBL_6_padClk;
wire CLK_int_0__CAND0_BLSBL_7_padClk;
wire CLK_int_0__CAND0_BLSBL_8_padClk;
wire CLK_int_0__CAND0_BLSBR_10_padClk;
wire CLK_int_0__CAND0_BLSBR_11_padClk;
wire CLK_int_0__CAND0_BLSBR_12_padClk;
wire CLK_int_0__CAND0_BLSBR_13_padClk;
wire CLK_int_0__CAND0_BLSBR_14_padClk;
wire CLK_int_0__CAND0_BLSBR_15_padClk;
wire CLK_int_0__CAND0_BLSBR_9_padClk;
wire CLK_int_0__CAND0_BLSTL_1_padClk;
wire CLK_int_0__CAND0_BLSTL_2_padClk;
wire CLK_int_0__CAND0_BLSTL_3_padClk;
wire CLK_int_0__CAND0_BLSTL_4_padClk;
wire CLK_int_0__CAND0_BLSTL_5_padClk;
wire CLK_int_0__CAND0_BLSTL_6_padClk;
wire CLK_int_0__CAND0_BLSTL_7_padClk;
wire CLK_int_0__CAND0_BLSTL_8_padClk;
wire CLK_int_0__CAND0_BLSTR_10_padClk;
wire CLK_int_0__CAND0_BLSTR_11_padClk;
wire CLK_int_0__CAND0_BLSTR_12_padClk;
wire CLK_int_0__CAND0_BLSTR_13_padClk;
wire CLK_int_0__CAND0_BLSTR_14_padClk;
wire CLK_int_0__CAND0_BLSTR_15_padClk;
wire CLK_int_0__CAND0_BLSTR_16_padClk;
wire CLK_int_0__CAND0_BLSTR_9_padClk;
wire CLK_int_0__CAND0_BRSBL_17_padClk;
wire CLK_int_0__CAND0_BRSBL_18_padClk;
wire CLK_int_0__CAND0_BRSBL_19_padClk;
wire CLK_int_0__CAND0_BRSBL_20_padClk;
wire CLK_int_0__CAND0_BRSBL_21_padClk;
wire CLK_int_0__CAND0_BRSBL_22_padClk;
wire CLK_int_0__CAND0_BRSBL_23_padClk;
wire CLK_int_0__CAND0_BRSBL_24_padClk;
wire CLK_int_0__CAND0_BRSBR_25_padClk;
wire CLK_int_0__CAND0_BRSBR_26_padClk;
wire CLK_int_0__CAND0_BRSBR_27_padClk;
wire CLK_int_0__CAND0_BRSBR_28_padClk;
wire CLK_int_0__CAND0_BRSBR_29_padClk;
wire CLK_int_0__CAND0_BRSTL_17_padClk;
wire CLK_int_0__CAND0_BRSTL_18_padClk;
wire CLK_int_0__CAND0_BRSTL_19_padClk;
wire CLK_int_0__CAND0_BRSTL_20_padClk;
wire CLK_int_0__CAND0_BRSTL_21_padClk;
wire CLK_int_0__CAND0_BRSTL_22_padClk;
wire CLK_int_0__CAND0_BRSTL_23_padClk;
wire CLK_int_0__CAND0_BRSTL_24_padClk;
wire CLK_int_0__CAND0_BRSTR_25_padClk;
wire CLK_int_0__CAND0_BRSTR_26_padClk;
wire CLK_int_0__CAND0_BRSTR_27_padClk;
wire CLK_int_0__CAND0_BRSTR_28_padClk;
wire CLK_int_0__CAND0_BRSTR_29_padClk;
wire CLK_int_0__CAND0_BRSTR_33_padClk;
wire CLK_int_0__CAND0_TLSBL_0_padClk;
wire CLK_int_0__CAND0_TLSBL_1_padClk;
wire CLK_int_0__CAND0_TLSBL_2_padClk;
wire CLK_int_0__CAND0_TLSBL_3_padClk;
wire CLK_int_0__CAND0_TLSBL_4_padClk;
wire CLK_int_0__CAND0_TLSBL_5_padClk;
wire CLK_int_0__CAND0_TLSBL_6_padClk;
wire CLK_int_0__CAND0_TLSBL_7_padClk;
wire CLK_int_0__CAND0_TLSBL_8_padClk;
wire CLK_int_0__CAND0_TLSBR_10_padClk;
wire CLK_int_0__CAND0_TLSBR_11_padClk;
wire CLK_int_0__CAND0_TLSBR_12_padClk;
wire CLK_int_0__CAND0_TLSBR_13_padClk;
wire CLK_int_0__CAND0_TLSBR_14_padClk;
wire CLK_int_0__CAND0_TLSBR_15_padClk;
wire CLK_int_0__CAND0_TLSBR_16_padClk;
wire CLK_int_0__CAND0_TLSBR_9_padClk;
wire CLK_int_0__CAND0_TLSTL_1_padClk;
wire CLK_int_0__CAND0_TLSTL_2_padClk;
wire CLK_int_0__CAND0_TLSTL_3_padClk;
wire CLK_int_0__CAND0_TLSTL_4_padClk;
wire CLK_int_0__CAND0_TLSTL_5_padClk;
wire CLK_int_0__CAND0_TLSTL_6_padClk;
wire CLK_int_0__CAND0_TLSTL_7_padClk;
wire CLK_int_0__CAND0_TLSTL_8_padClk;
wire CLK_int_0__CAND0_TLSTR_10_padClk;
wire CLK_int_0__CAND0_TLSTR_11_padClk;
wire CLK_int_0__CAND0_TLSTR_12_padClk;
wire CLK_int_0__CAND0_TLSTR_13_padClk;
wire CLK_int_0__CAND0_TLSTR_14_padClk;
wire CLK_int_0__CAND0_TLSTR_15_padClk;
wire CLK_int_0__CAND0_TLSTR_16_padClk;
wire CLK_int_0__CAND0_TLSTR_9_padClk;
wire CLK_int_0__CAND0_TRSBL_17_padClk;
wire CLK_int_0__CAND0_TRSBL_18_padClk;
wire CLK_int_0__CAND0_TRSBL_19_padClk;
wire CLK_int_0__CAND0_TRSBL_21_padClk;
wire CLK_int_0__CAND0_TRSBL_22_padClk;
wire CLK_int_0__CAND0_TRSBL_23_padClk;
wire CLK_int_0__CAND0_TRSBL_24_padClk;
wire CLK_int_0__CAND0_TRSBR_25_padClk;
wire CLK_int_0__CAND0_TRSBR_26_padClk;
wire CLK_int_0__CAND0_TRSBR_27_padClk;
wire CLK_int_0__CAND0_TRSBR_28_padClk;
wire CLK_int_0__CAND0_TRSBR_29_padClk;
wire CLK_int_0__CAND0_TRSBR_33_padClk;
wire CLK_int_0__CAND0_TRSTL_17_padClk;
wire CLK_int_0__CAND0_TRSTL_18_padClk;
wire CLK_int_0__CAND0_TRSTL_19_padClk;
wire CLK_int_0__CAND0_TRSTL_20_padClk;
wire CLK_int_0__CAND0_TRSTL_21_padClk;
wire CLK_int_0__CAND0_TRSTL_22_padClk;
wire CLK_int_0__CAND0_TRSTL_23_padClk;
wire CLK_int_0__CAND0_TRSTL_24_padClk;
wire CLK_int_0__CAND0_TRSTR_25_padClk;
wire CLK_int_0__CAND0_TRSTR_26_padClk;
wire CLK_int_0__CAND0_TRSTR_27_padClk;
wire CLK_int_0__CAND0_TRSTR_28_padClk;
wire CLK_int_0__CAND0_TRSTR_29_padClk;
wire CLK_int_0__CAND0_TRSTR_33_padClk;
wire CLK_int_0__GMUX_0_padClk;
wire CLK_int_0__QMUX_BL0_padClk;
wire CLK_int_0__QMUX_BR0_padClk;
wire CLK_int_0__QMUX_TL0_padClk;
wire CLK_int_0__QMUX_TR0_padClk;
wire CLK_int_0__SQMUX_BLSBL0_padClk;
wire CLK_int_0__SQMUX_BLSBR0_padClk;
wire CLK_int_0__SQMUX_BLSTL0_padClk;
wire CLK_int_0__SQMUX_BLSTR0_padClk;
wire CLK_int_0__SQMUX_BRSBL0_padClk;
wire CLK_int_0__SQMUX_BRSBR0_padClk;
wire CLK_int_0__SQMUX_BRSTL0_padClk;
wire CLK_int_0__SQMUX_BRSTR0_padClk;
wire CLK_int_0__SQMUX_TLSBL0_padClk;
wire CLK_int_0__SQMUX_TLSBR0_padClk;
wire CLK_int_0__SQMUX_TLSTL0_padClk;
wire CLK_int_0__SQMUX_TLSTR0_padClk;
wire CLK_int_0__SQMUX_TRSBL0_padClk;
wire CLK_int_0__SQMUX_TRSBR0_padClk;
wire CLK_int_0__SQMUX_TRSTL0_padClk;
wire CLK_int_0__SQMUX_TRSTR0_padClk;
wire CLK_int_1__CAND1_BRSTL_20_padClk;
wire CLK_int_1__CAND1_BRSTL_21_padClk;
wire CLK_int_1__GMUX_1_padClk;
wire CLK_int_1__QMUX_BR1_padClk;
wire CLK_int_1__SQMUX_BRSTL1_padClk;
wire CLK_int_2__CAND2_TRSBL_18_padClk;
wire CLK_int_2__GMUX_2_padClk;
wire CLK_int_2__QMUX_TR2_padClk;
wire CLK_int_2__SQMUX_TRSBL2_padClk;
wire CLK_int_3__CAND3_TRSBL_17_padClk;
wire CLK_int_3__GMUX_3_padClk;
wire CLK_int_3__QMUX_TR3_padClk;
wire CLK_int_3__SQMUX_TRSBL3_padClk;
wire CLK_int_4__CAND4_TRSBL_20_padClk;
wire CLK_int_4__GMUX_4_padClk;
wire CLK_int_4__QMUX_TR4_padClk;
wire CLK_int_4__SQMUX_TRSBL4_padClk;
wire CLK_int_5__CAND5_TRSBL_17_padClk;
wire CLK_int_5__GMUX_5_padClk;
wire CLK_int_5__QMUX_TR5_padClk;
wire CLK_int_5__SQMUX_TRSBL5_padClk;
wire NET_0;
wire NET_0_CAND1_BRSBR_25_tpGCLKBUF;
wire NET_0_CAND1_BRSBR_26_tpGCLKBUF;
wire NET_0_CAND1_BRSBR_27_tpGCLKBUF;
wire NET_0_CAND1_BRSBR_28_tpGCLKBUF;
wire NET_0_CAND1_BRSBR_29_tpGCLKBUF;
wire NET_0_SQMUX_BRSBR1_tpGCLKBUF;
wire NET_1;
wire NET_10;
wire NET_100;
wire NET_101;
wire NET_102;
wire NET_103;
wire NET_104;
wire NET_105;
wire NET_106;
wire NET_107;
wire NET_108;
wire NET_109;
wire NET_11;
wire NET_110;
wire NET_111;
wire NET_112;
wire NET_113;
wire NET_113_CAND4_BRSBL_17_tpGCLKBUF;
wire NET_113_CAND4_BRSBL_18_tpGCLKBUF;
wire NET_113_CAND4_BRSBL_19_tpGCLKBUF;
wire NET_113_CAND4_BRSBL_20_tpGCLKBUF;
wire NET_113_SQMUX_BRSBL4_tpGCLKBUF;
wire NET_114;
wire NET_115;
wire NET_116;
wire NET_117;
wire NET_118;
wire NET_119;
wire NET_12;
wire NET_120;
wire NET_121;
wire NET_122;
wire NET_123;
wire NET_124;
wire NET_125;
wire NET_126;
wire NET_126_CAND3_TLSBR_10_tpGCLKBUF;
wire NET_126_CAND3_TLSBR_11_tpGCLKBUF;
wire NET_126_CAND3_TLSBR_12_tpGCLKBUF;
wire NET_126_CAND3_TLSBR_13_tpGCLKBUF;
wire NET_126_CAND3_TLSBR_14_tpGCLKBUF;
wire NET_126_SQMUX_TLSBR3_tpGCLKBUF;
wire NET_127;
wire NET_127_CAND4_TLSBR_10_tpGCLKBUF;
wire NET_127_CAND4_TLSBR_12_tpGCLKBUF;
wire NET_127_CAND4_TLSBR_13_tpGCLKBUF;
wire NET_127_CAND4_TLSBR_14_tpGCLKBUF;
wire NET_127_CAND4_TLSBR_15_tpGCLKBUF;
wire NET_127_CAND4_TLSBR_9_tpGCLKBUF;
wire NET_127_SQMUX_TLSBR4_tpGCLKBUF;
wire NET_128;
wire NET_129;
wire NET_13;
wire NET_130;
wire NET_131;
wire NET_132;
wire NET_133;
wire NET_134;
wire NET_135;
wire NET_136;
wire NET_137;
wire NET_138;
wire NET_139;
wire NET_14;
wire NET_140;
wire NET_141;
wire NET_142;
wire NET_143;
wire NET_144;
wire NET_145;
wire NET_146;
wire NET_147;
wire NET_148;
wire NET_149;
wire NET_15;
wire NET_150;
wire NET_151;
wire NET_152;
wire NET_153;
wire NET_154;
wire NET_155;
wire NET_156;
wire NET_157;
wire NET_158;
wire NET_159;
wire NET_16;
wire NET_160;
wire NET_161;
wire NET_162;
wire NET_163;
wire NET_164;
wire NET_165;
wire NET_166;
wire NET_167;
wire NET_168;
wire NET_169;
wire NET_17;
wire NET_170;
wire NET_171;
wire NET_172;
wire NET_173;
wire NET_174;
wire NET_175;
wire NET_176;
wire NET_177;
wire NET_178;
wire NET_179;
wire NET_18;
wire NET_180;
wire NET_181;
wire NET_182;
wire NET_183;
wire NET_184;
wire NET_185;
wire NET_186;
wire NET_187;
wire NET_188;
wire NET_189;
wire NET_19;
wire NET_190;
wire NET_191;
wire NET_192;
wire NET_193;
wire NET_194;
wire NET_195;
wire NET_196;
wire NET_197;
wire NET_198;
wire NET_199;
wire NET_2;
wire NET_20;
wire NET_200;
wire NET_201;
wire NET_202;
wire NET_203;
wire NET_204;
wire NET_205;
wire NET_206;
wire NET_207;
wire NET_208;
wire NET_209;
wire NET_21;
wire NET_210;
wire NET_211;
wire NET_212;
wire NET_213;
wire NET_214;
wire NET_215;
wire NET_216;
wire NET_217;
wire NET_218;
wire NET_219;
wire NET_21_CAND4_BLSTR_12_tpGCLKBUF;
wire NET_21_CAND4_BLSTR_13_tpGCLKBUF;
wire NET_21_CAND4_BLSTR_15_tpGCLKBUF;
wire NET_21_SQMUX_BLSTR4_tpGCLKBUF;
wire NET_22;
wire NET_220;
wire NET_221;
wire NET_222;
wire NET_223;
wire NET_224;
wire NET_225;
wire NET_226;
wire NET_227;
wire NET_228;
wire NET_229;
wire NET_23;
wire NET_230;
wire NET_231;
wire NET_232;
wire NET_233;
wire NET_234;
wire NET_235;
wire NET_236;
wire NET_237;
wire NET_238;
wire NET_239;
wire NET_24;
wire NET_240;
wire NET_241;
wire NET_242;
wire NET_243;
wire NET_244;
wire NET_245;
wire NET_246;
wire NET_247;
wire NET_248;
wire NET_249;
wire NET_25;
wire NET_250;
wire NET_251;
wire NET_252;
wire NET_253;
wire NET_254;
wire NET_255;
wire NET_256;
wire NET_257;
wire NET_258;
wire NET_259;
wire NET_26;
wire NET_260;
wire NET_261;
wire NET_262;
wire NET_263;
wire NET_264;
wire NET_265;
wire NET_266;
wire NET_267;
wire NET_268;
wire NET_269;
wire NET_27;
wire NET_270;
wire NET_271;
wire NET_272;
wire NET_273;
wire NET_274;
wire NET_275;
wire NET_276;
wire NET_277;
wire NET_278;
wire NET_279;
wire NET_27_CAND5_BLSTR_10_tpGCLKBUF;
wire NET_27_CAND5_BLSTR_11_tpGCLKBUF;
wire NET_27_CAND5_BLSTR_12_tpGCLKBUF;
wire NET_27_CAND5_BLSTR_14_tpGCLKBUF;
wire NET_27_CAND5_BLSTR_15_tpGCLKBUF;
wire NET_27_SQMUX_BLSTR5_tpGCLKBUF;
wire NET_28;
wire NET_280;
wire NET_281;
wire NET_282;
wire NET_283;
wire NET_284;
wire NET_285;
wire NET_286;
wire NET_287;
wire NET_288;
wire NET_289;
wire NET_29;
wire NET_290;
wire NET_291;
wire NET_292;
wire NET_293;
wire NET_294;
wire NET_295;
wire NET_296;
wire NET_297;
wire NET_298;
wire NET_299;
wire NET_3;
wire NET_30;
wire NET_300;
wire NET_301;
wire NET_302;
wire NET_303;
wire NET_304;
wire NET_305;
wire NET_306;
wire NET_307;
wire NET_308;
wire NET_309;
wire NET_30_CAND5_TLSBR_10_tpGCLKBUF;
wire NET_30_CAND5_TLSBR_11_tpGCLKBUF;
wire NET_30_SQMUX_TLSBR5_tpGCLKBUF;
wire NET_31;
wire NET_310;
wire NET_311;
wire NET_312;
wire NET_313;
wire NET_314;
wire NET_315;
wire NET_316;
wire NET_317;
wire NET_318;
wire NET_319;
wire NET_32;
wire NET_320;
wire NET_321;
wire NET_322;
wire NET_323;
wire NET_324;
wire NET_325;
wire NET_326;
wire NET_327;
wire NET_328;
wire NET_329;
wire NET_33;
wire NET_330;
wire NET_331;
wire NET_332;
wire NET_333;
wire NET_334;
wire NET_335;
wire NET_336;
wire NET_337;
wire NET_338;
wire NET_339;
wire NET_33_CAND2_TLSBR_10_tpGCLKBUF;
wire NET_33_CAND2_TLSBR_11_tpGCLKBUF;
wire NET_33_CAND2_TLSBR_12_tpGCLKBUF;
wire NET_33_CAND2_TLSBR_14_tpGCLKBUF;
wire NET_33_CAND2_TLSBR_16_tpGCLKBUF;
wire NET_33_SQMUX_TLSBR2_tpGCLKBUF;
wire NET_34;
wire NET_340;
wire NET_341;
wire NET_342;
wire NET_343;
wire NET_344;
wire NET_345;
wire NET_346;
wire NET_347;
wire NET_348;
wire NET_349;
wire NET_35;
wire NET_350;
wire NET_351;
wire NET_352;
wire NET_353;
wire NET_354;
wire NET_355;
wire NET_356;
wire NET_357;
wire NET_358;
wire NET_359;
wire NET_36;
wire NET_360;
wire NET_361;
wire NET_362;
wire NET_363;
wire NET_364;
wire NET_365;
wire NET_366;
wire NET_367;
wire NET_368;
wire NET_369;
wire NET_37;
wire NET_370;
wire NET_371;
wire NET_372;
wire NET_373;
wire NET_374;
wire NET_375;
wire NET_376;
wire NET_377;
wire NET_378;
wire NET_379;
wire NET_38;
wire NET_380;
wire NET_381;
wire NET_382;
wire NET_383;
wire NET_384;
wire NET_385;
wire NET_386;
wire NET_387;
wire NET_388;
wire NET_389;
wire NET_39;
wire NET_390;
wire NET_391;
wire NET_392;
wire NET_393;
wire NET_394;
wire NET_395;
wire NET_396;
wire NET_397;
wire NET_398;
wire NET_399;
wire NET_4;
wire NET_40;
wire NET_400;
wire NET_401;
wire NET_402;
wire NET_403;
wire NET_404;
wire NET_405;
wire NET_406;
wire NET_407;
wire NET_408;
wire NET_409;
wire NET_41;
wire NET_410;
wire NET_411;
wire NET_412;
wire NET_413;
wire NET_414;
wire NET_415;
wire NET_416;
wire NET_417;
wire NET_418;
wire NET_419;
wire NET_42;
wire NET_420;
wire NET_421;
wire NET_422;
wire NET_423;
wire NET_424;
wire NET_425;
wire NET_426;
wire NET_427;
wire NET_428;
wire NET_429;
wire NET_43;
wire NET_430;
wire NET_431;
wire NET_432;
wire NET_433;
wire NET_434;
wire NET_435;
wire NET_436;
wire NET_437;
wire NET_438;
wire NET_439;
wire NET_44;
wire NET_440;
wire NET_441;
wire NET_442;
wire NET_443;
wire NET_444;
wire NET_445;
wire NET_446;
wire NET_447;
wire NET_448;
wire NET_449;
wire NET_45;
wire NET_450;
wire NET_451;
wire NET_452;
wire NET_453;
wire NET_454;
wire NET_455;
wire NET_456;
wire NET_457;
wire NET_458;
wire NET_459;
wire NET_46;
wire NET_460;
wire NET_461;
wire NET_462;
wire NET_463;
wire NET_464;
wire NET_465;
wire NET_466;
wire NET_467;
wire NET_468;
wire NET_469;
wire NET_47;
wire NET_470;
wire NET_471;
wire NET_472;
wire NET_473;
wire NET_474;
wire NET_475;
wire NET_476;
wire NET_477;
wire NET_478;
wire NET_479;
wire NET_48;
wire NET_480;
wire NET_481;
wire NET_482;
wire NET_482_CAND3_BLSBL_5_tpGCLKBUF;
wire NET_482_CAND3_BLSBL_6_tpGCLKBUF;
wire NET_482_CAND3_BLSBL_8_tpGCLKBUF;
wire NET_482_SQMUX_BLSBL3_tpGCLKBUF;
wire NET_483;
wire NET_484;
wire NET_485;
wire NET_486;
wire NET_487;
wire NET_488;
wire NET_489;
wire NET_49;
wire NET_490;
wire NET_491;
wire NET_492;
wire NET_493;
wire NET_494;
wire NET_495;
wire NET_496;
wire NET_497;
wire NET_498;
wire NET_499;
wire NET_5;
wire NET_50;
wire NET_500;
wire NET_501;
wire NET_502;
wire NET_503;
wire NET_504;
wire NET_505;
wire NET_506;
wire NET_507;
wire NET_508;
wire NET_509;
wire NET_51;
wire NET_510;
wire NET_511;
wire NET_512;
wire NET_513;
wire NET_514;
wire NET_515;
wire NET_516;
wire NET_517;
wire NET_518;
wire NET_519;
wire NET_52;
wire NET_520;
wire NET_521;
wire NET_522;
wire NET_523;
wire NET_524;
wire NET_525;
wire NET_526;
wire NET_527;
wire NET_528;
wire NET_529;
wire NET_53;
wire NET_530;
wire NET_531;
wire NET_532;
wire NET_533;
wire NET_534;
wire NET_535;
wire NET_536;
wire NET_537;
wire NET_538;
wire NET_539;
wire NET_54;
wire NET_540;
wire NET_541;
wire NET_542;
wire NET_543;
wire NET_544;
wire NET_545;
wire NET_546;
wire NET_547;
wire NET_548;
wire NET_549;
wire NET_55;
wire NET_550;
wire NET_551;
wire NET_552;
wire NET_553;
wire NET_554;
wire NET_555;
wire NET_556;
wire NET_557;
wire NET_558;
wire NET_559;
wire NET_56;
wire NET_560;
wire NET_561;
wire NET_562;
wire NET_563;
wire NET_564;
wire NET_565;
wire NET_566;
wire NET_567;
wire NET_568;
wire NET_569;
wire NET_57;
wire NET_570;
wire NET_571;
wire NET_572;
wire NET_573;
wire NET_574;
wire NET_575;
wire NET_576;
wire NET_577;
wire NET_578;
wire NET_579;
wire NET_58;
wire NET_580;
wire NET_581;
wire NET_582;
wire NET_583;
wire NET_584;
wire NET_585;
wire NET_586;
wire NET_587;
wire NET_588;
wire NET_589;
wire NET_59;
wire NET_590;
wire NET_591;
wire NET_592;
wire NET_593;
wire NET_594;
wire NET_595;
wire NET_596;
wire NET_597;
wire NET_598;
wire NET_599;
wire NET_59_CAND5_TRSTL_19_tpGCLKBUF;
wire NET_59_CAND5_TRSTL_20_tpGCLKBUF;
wire NET_59_CAND5_TRSTL_21_tpGCLKBUF;
wire NET_59_SQMUX_TRSTL5_tpGCLKBUF;
wire NET_6;
wire NET_60;
wire NET_600;
wire NET_601;
wire NET_602;
wire NET_603;
wire NET_604;
wire NET_605;
wire NET_606;
wire NET_607;
wire NET_608;
wire NET_609;
wire NET_61;
wire NET_610;
wire NET_611;
wire NET_612;
wire NET_613;
wire NET_614;
wire NET_615;
wire NET_616;
wire NET_617;
wire NET_618;
wire NET_619;
wire NET_62;
wire NET_620;
wire NET_621;
wire NET_622;
wire NET_623;
wire NET_624;
wire NET_625;
wire NET_626;
wire NET_627;
wire NET_628;
wire NET_629;
wire NET_62_CAND3_BRSTL_17_tpGCLKBUF;
wire NET_62_CAND3_BRSTL_18_tpGCLKBUF;
wire NET_62_CAND3_BRSTL_19_tpGCLKBUF;
wire NET_62_CAND3_BRSTL_20_tpGCLKBUF;
wire NET_62_CAND3_BRSTL_21_tpGCLKBUF;
wire NET_62_SQMUX_BRSTL3_tpGCLKBUF;
wire NET_63;
wire NET_630;
wire NET_631;
wire NET_632;
wire NET_633;
wire NET_634;
wire NET_635;
wire NET_636;
wire NET_637;
wire NET_638;
wire NET_639;
wire NET_64;
wire NET_640;
wire NET_641;
wire NET_642;
wire NET_643;
wire NET_644;
wire NET_645;
wire NET_646;
wire NET_647;
wire NET_648;
wire NET_649;
wire NET_65;
wire NET_650;
wire NET_651;
wire NET_652;
wire NET_653;
wire NET_654;
wire NET_655;
wire NET_656;
wire NET_657;
wire NET_658;
wire NET_659;
wire NET_66;
wire NET_660;
wire NET_661;
wire NET_662;
wire NET_663;
wire NET_664;
wire NET_665;
wire NET_666;
wire NET_667;
wire NET_668;
wire NET_669;
wire NET_67;
wire NET_670;
wire NET_671;
wire NET_672;
wire NET_673;
wire NET_674;
wire NET_675;
wire NET_676;
wire NET_677;
wire NET_678;
wire NET_679;
wire NET_68;
wire NET_680;
wire NET_681;
wire NET_682;
wire NET_683;
wire NET_684;
wire NET_685;
wire NET_686;
wire NET_687;
wire NET_688;
wire NET_689;
wire NET_69;
wire NET_690;
wire NET_691;
wire NET_692;
wire NET_693;
wire NET_694;
wire NET_695;
wire NET_696;
wire NET_697;
wire NET_698;
wire NET_699;
wire NET_7;
wire NET_70;
wire NET_700;
wire NET_701;
wire NET_702;
wire NET_703;
wire NET_704;
wire NET_705;
wire NET_706;
wire NET_707;
wire NET_708;
wire NET_709;
wire NET_71;
wire NET_710;
wire NET_711;
wire NET_712;
wire NET_713;
wire NET_714;
wire NET_715;
wire NET_716;
wire NET_717;
wire NET_718;
wire NET_719;
wire NET_72;
wire NET_720;
wire NET_721;
wire NET_722;
wire NET_723;
wire NET_724;
wire NET_725;
wire NET_726;
wire NET_727;
wire NET_728;
wire NET_729;
wire NET_73;
wire NET_730;
wire NET_731;
wire NET_732;
wire NET_733;
wire NET_734;
wire NET_735;
wire NET_736;
wire NET_737;
wire NET_738;
wire NET_739;
wire NET_73_CAND3_TLSBL_1_tpGCLKBUF;
wire NET_73_CAND3_TLSBL_2_tpGCLKBUF;
wire NET_73_CAND3_TLSBL_3_tpGCLKBUF;
wire NET_73_CAND3_TLSBL_4_tpGCLKBUF;
wire NET_73_SQMUX_TLSBL3_tpGCLKBUF;
wire NET_74;
wire NET_740;
wire NET_741;
wire NET_742;
wire NET_743;
wire NET_744;
wire NET_745;
wire NET_746;
wire NET_747;
wire NET_748;
wire NET_749;
wire NET_75;
wire NET_750;
wire NET_751;
wire NET_752;
wire NET_753;
wire NET_754;
wire NET_755;
wire NET_756;
wire NET_757;
wire NET_758;
wire NET_759;
wire NET_75_CAND5_TLSBL_1_tpGCLKBUF;
wire NET_75_CAND5_TLSBL_2_tpGCLKBUF;
wire NET_75_CAND5_TLSBL_3_tpGCLKBUF;
wire NET_75_CAND5_TLSBL_6_tpGCLKBUF;
wire NET_75_SQMUX_TLSBL5_tpGCLKBUF;
wire NET_76;
wire NET_760;
wire NET_761;
wire NET_762;
wire NET_763;
wire NET_764;
wire NET_765;
wire NET_766;
wire NET_767;
wire NET_768;
wire NET_769;
wire NET_77;
wire NET_770;
wire NET_771;
wire NET_772;
wire NET_773;
wire NET_774;
wire NET_775;
wire NET_776;
wire NET_777;
wire NET_778;
wire NET_779;
wire NET_78;
wire NET_780;
wire NET_781;
wire NET_782;
wire NET_783;
wire NET_784;
wire NET_785;
wire NET_786;
wire NET_787;
wire NET_788;
wire NET_789;
wire NET_79;
wire NET_790;
wire NET_791;
wire NET_792;
wire NET_793;
wire NET_794;
wire NET_795;
wire NET_796;
wire NET_797;
wire NET_798;
wire NET_799;
wire NET_8;
wire NET_80;
wire NET_800;
wire NET_801;
wire NET_802;
wire NET_803;
wire NET_804;
wire NET_805;
wire NET_806;
wire NET_807;
wire NET_808;
wire NET_809;
wire NET_81;
wire NET_810;
wire NET_811;
wire NET_812;
wire NET_813;
wire NET_814;
wire NET_815;
wire NET_816;
wire NET_817;
wire NET_818;
wire NET_819;
wire NET_82;
wire NET_820;
wire NET_821;
wire NET_822;
wire NET_823;
wire NET_824;
wire NET_825;
wire NET_826;
wire NET_827;
wire NET_828;
wire NET_829;
wire NET_83;
wire NET_830;
wire NET_831;
wire NET_832;
wire NET_833;
wire NET_834;
wire NET_835;
wire NET_836;
wire NET_837;
wire NET_838;
wire NET_839;
wire NET_84;
wire NET_840;
wire NET_841;
wire NET_842;
wire NET_843;
wire NET_844;
wire NET_845;
wire NET_846;
wire NET_847;
wire NET_848;
wire NET_849;
wire NET_85;
wire NET_850;
wire NET_851;
wire NET_852;
wire NET_853;
wire NET_854;
wire NET_855;
wire NET_856;
wire NET_857;
wire NET_858;
wire NET_859;
wire NET_86;
wire NET_860;
wire NET_861;
wire NET_862;
wire NET_863;
wire NET_864;
wire NET_865;
wire NET_866;
wire NET_867;
wire NET_868;
wire NET_869;
wire NET_87;
wire NET_870;
wire NET_871;
wire NET_872;
wire NET_873;
wire NET_874;
wire NET_875;
wire NET_876;
wire NET_877;
wire NET_878;
wire NET_879;
wire NET_88;
wire NET_880;
wire NET_881;
wire NET_882;
wire NET_883;
wire NET_884;
wire NET_885;
wire NET_886;
wire NET_887;
wire NET_888;
wire NET_889;
wire NET_89;
wire NET_890;
wire NET_891;
wire NET_892;
wire NET_893;
wire NET_894;
wire NET_895;
wire NET_896;
wire NET_897;
wire NET_898;
wire NET_899;
wire NET_9;
wire NET_90;
wire NET_900;
wire NET_901;
wire NET_902;
wire NET_903;
wire NET_904;
wire NET_905;
wire NET_906;
wire NET_907;
wire NET_908;
wire NET_909;
wire NET_91;
wire NET_910;
wire NET_911;
wire NET_912;
wire NET_913;
wire NET_914;
wire NET_915;
wire NET_916;
wire NET_917;
wire NET_918;
wire NET_919;
wire NET_92;
wire NET_920;
wire NET_921;
wire NET_922;
wire NET_923;
wire NET_924;
wire NET_925;
wire NET_926;
wire NET_927;
wire NET_928;
wire NET_929;
wire NET_93;
wire NET_930;
wire NET_94;
wire NET_95;
wire NET_96;
wire NET_97;
wire NET_98;
wire NET_99;
wire apb_fsm_0__CAND4_BRSTL_17_tpGCLKBUF;
wire apb_fsm_0__CAND4_BRSTL_18_tpGCLKBUF;
wire apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF;
wire apb_fsm_0__CAND4_BRSTL_20_tpGCLKBUF;
wire apb_fsm_0__SQMUX_BRSTL4_tpGCLKBUF;
wire launch_p0;
wire launch_p1;
wire launch_p2;
wire launch_p3;
wire lint_ADDR_int_11__CAND4_TLSBL_1_tpGCLKBUF;
wire lint_ADDR_int_11__CAND4_TLSBL_2_tpGCLKBUF;
wire lint_ADDR_int_11__CAND4_TLSBL_6_tpGCLKBUF;
wire lint_ADDR_int_11__SQMUX_TLSBL4_tpGCLKBUF;
wire lint_ADDR_int_13__CAND5_BRSTL_18_tpGCLKBUF;
wire lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF;
wire lint_ADDR_int_13__CAND5_BRSTL_20_tpGCLKBUF;
wire lint_ADDR_int_13__SQMUX_BRSTL5_tpGCLKBUF;
wire lint_ADDR_int_2__CAND3_BLSTR_11_tpGCLKBUF;
wire lint_ADDR_int_2__CAND3_BLSTR_12_tpGCLKBUF;
wire lint_ADDR_int_2__CAND3_BLSTR_14_tpGCLKBUF;
wire lint_ADDR_int_2__CAND3_BLSTR_15_tpGCLKBUF;
wire lint_ADDR_int_2__CAND3_BLSTR_16_tpGCLKBUF;
wire lint_ADDR_int_2__SQMUX_BLSTR3_tpGCLKBUF;
wire lint_GNT;
wire lint_GNT_dup_0;
wire lint_REQ;
wire lint_REQ_int;
wire lint_VALID;
wire lint_VALID_dup_0;
wire lint_WEN;
wire lint_WEN_int;
wire lint_clk;
wire m0_coef_powerdn;
wire m0_coef_rclk;
wire m0_coef_wclk;
wire m0_coef_wdsel;
wire m0_coef_wdsel_dup_0;
wire m0_coef_we;
wire m0_coef_we_dup_0;
wire m0_m0_clk;
wire m0_m0_clken;
wire m0_m0_clken_dup_0;
wire m0_m0_clr;
wire m0_m0_clr_dup_0;
wire m0_m0_csel;
wire m0_m0_csel_dup_0;
wire m0_m0_osel;
wire m0_m0_osel_dup_0;
wire m0_m0_reset;
wire m0_m0_reset_dup_0;
wire m0_m0_rnd;
wire m0_m0_rnd_dup_0;
wire m0_m0_sat;
wire m0_m0_sat_dup_0;
wire m0_m0_tc;
wire m0_m0_tc_dup_0;
wire m0_m1_clk;
wire m0_m1_clken;
wire m0_m1_clken_dup_0;
wire m0_m1_clr;
wire m0_m1_clr_dup_0;
wire m0_m1_csel;
wire m0_m1_csel_dup_0;
wire m0_m1_osel;
wire m0_m1_osel_dup_0;
wire m0_m1_reset;
wire m0_m1_reset_dup_0;
wire m0_m1_rnd;
wire m0_m1_rnd_dup_0;
wire m0_m1_sat;
wire m0_m1_sat_dup_0;
wire m0_m1_tc;
wire m0_m1_tc_dup_0;
wire m0_oper0_powerdn;
wire m0_oper0_rclk;
wire m0_oper0_wclk;
wire m0_oper0_wdsel;
wire m0_oper0_wdsel_dup_0;
wire m0_oper0_we;
wire m0_oper0_we_dup_0;
wire m0_oper1_powerdn;
wire m0_oper1_rclk;
wire m0_oper1_wclk;
wire m0_oper1_wdsel;
wire m0_oper1_wdsel_dup_0;
wire m0_oper1_we;
wire m0_oper1_we_dup_0;
wire m1_coef_powerdn;
wire m1_coef_rclk;
wire m1_coef_wclk;
wire m1_coef_wdsel;
wire m1_coef_wdsel_dup_0;
wire m1_coef_we;
wire m1_coef_we_dup_0;
wire m1_m0_clk;
wire m1_m0_clken;
wire m1_m0_clken_dup_0;
wire m1_m0_clr;
wire m1_m0_clr_dup_0;
wire m1_m0_csel;
wire m1_m0_csel_dup_0;
wire m1_m0_osel;
wire m1_m0_osel_dup_0;
wire m1_m0_reset;
wire m1_m0_reset_dup_0;
wire m1_m0_rnd;
wire m1_m0_rnd_dup_0;
wire m1_m0_sat;
wire m1_m0_sat_dup_0;
wire m1_m0_tc;
wire m1_m0_tc_dup_0;
wire m1_m1_clk;
wire m1_m1_clken;
wire m1_m1_clken_dup_0;
wire m1_m1_clr;
wire m1_m1_clr_dup_0;
wire m1_m1_csel;
wire m1_m1_csel_dup_0;
wire m1_m1_osel;
wire m1_m1_osel_dup_0;
wire m1_m1_reset;
wire m1_m1_reset_dup_0;
wire m1_m1_rnd;
wire m1_m1_rnd_dup_0;
wire m1_m1_sat;
wire m1_m1_sat_dup_0;
wire m1_m1_tc;
wire m1_m1_tc_dup_0;
wire m1_oper0_powerdn;
wire m1_oper0_rclk;
wire m1_oper0_wclk;
wire m1_oper0_wdsel;
wire m1_oper0_wdsel_dup_0;
wire m1_oper0_we;
wire m1_oper0_we_dup_0;
wire m1_oper1_powerdn;
wire m1_oper1_rclk;
wire m1_oper1_wclk;
wire m1_oper1_wdsel;
wire m1_oper1_wdsel_dup_0;
wire m1_oper1_we;
wire m1_oper1_we_dup_0;
wire not_RESET_0;
wire not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF;
wire not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF;
wire not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_22_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF;
wire not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBL_17_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBL_18_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBL_19_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBL_20_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBR_27_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBR_28_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSBR_29_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTL_21_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF;
wire not_RESET_0_CAND2_BRSTR_29_tpGCLKBUF;
wire not_RESET_0_QMUX_BL1_tpGCLKBUF;
wire not_RESET_0_QMUX_BR2_tpGCLKBUF;
wire not_RESET_0_QMUX_TL1_tpGCLKBUF;
wire not_RESET_0_QMUX_TR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSBL2_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSBR2_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSTL2_tpGCLKBUF;
wire not_RESET_0_SQMUX_BRSTR2_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSBL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF;
wire not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF;
wire not_RESET_1;
wire not_RESET_2;
wire not_RESET_3;
wire not_apb_fsm_0;
wire not_apb_fsm_1;
wire not_p3_fsm_0;
wire not_tcdm_wen_p0;
wire not_tcdm_wen_p1;
wire not_tcdm_wen_p2;
wire nx10146z1;
wire nx10146z2;
wire nx10406z1;
wire nx10775z1;
wire nx11310z3;
wire nx11311z1;
wire nx11311z1_CAND5_BRSBL_17_tpGCLKBUF;
wire nx11311z1_CAND5_BRSBL_18_tpGCLKBUF;
wire nx11311z1_CAND5_BRSBL_19_tpGCLKBUF;
wire nx11311z1_CAND5_BRSBL_20_tpGCLKBUF;
wire nx11311z1_SQMUX_BRSBL5_tpGCLKBUF;
wire nx11311z2;
wire nx11311z3;
wire nx11312z1;
wire nx11312z1_CAND3_TRSTR_25_tpGCLKBUF;
wire nx11312z1_CAND3_TRSTR_26_tpGCLKBUF;
wire nx11312z1_CAND3_TRSTR_27_tpGCLKBUF;
wire nx11312z1_CAND3_TRSTR_28_tpGCLKBUF;
wire nx11312z1_CAND3_TRSTR_29_tpGCLKBUF;
wire nx11312z1_CAND4_TRSBR_25_tpGCLKBUF;
wire nx11312z1_CAND4_TRSBR_26_tpGCLKBUF;
wire nx11312z1_CAND4_TRSBR_27_tpGCLKBUF;
wire nx11312z1_CAND4_TRSBR_28_tpGCLKBUF;
wire nx11312z1_CAND4_TRSBR_29_tpGCLKBUF;
wire nx11312z1_SQMUX_TRSBR4_tpGCLKBUF;
wire nx11312z1_SQMUX_TRSTR3_tpGCLKBUF;
wire nx11312z3;
wire nx11312z5;
wire nx11313z1;
wire nx11313z1_CAND2_TRSTL_17_tpGCLKBUF;
wire nx11313z1_CAND2_TRSTL_18_tpGCLKBUF;
wire nx11313z1_CAND2_TRSTL_19_tpGCLKBUF;
wire nx11313z1_CAND2_TRSTL_20_tpGCLKBUF;
wire nx11313z1_CAND2_TRSTL_21_tpGCLKBUF;
wire nx11313z1_SQMUX_TRSTL2_tpGCLKBUF;
wire nx11313z3;
wire nx11313z5;
wire nx12574z1;
wire nx12783z2;
wire nx12783z2_CAND4_BLSTL_5_tpGCLKBUF;
wire nx12783z2_CAND4_BLSTL_6_tpGCLKBUF;
wire nx12783z2_CAND4_BLSTL_7_tpGCLKBUF;
wire nx12783z2_CAND4_BLSTL_8_tpGCLKBUF;
wire nx12783z2_SQMUX_BLSTL4_tpGCLKBUF;
wire nx12973z2;
wire nx12973z2_CAND3_TRSBR_26_tpGCLKBUF;
wire nx12973z2_CAND3_TRSBR_27_tpGCLKBUF;
wire nx12973z2_SQMUX_TRSBR3_tpGCLKBUF;
wire nx13379z2;
wire nx13970z2;
wire nx13970z2_CAND2_TRSBR_26_tpGCLKBUF;
wire nx13970z2_CAND2_TRSBR_27_tpGCLKBUF;
wire nx13970z2_CAND2_TRSBR_28_tpGCLKBUF;
wire nx13970z2_SQMUX_TRSBR2_tpGCLKBUF;
wire nx14650z1;
wire nx14650z1_CAND3_BLSBR_14_tpGCLKBUF;
wire nx14650z1_CAND3_BLSBR_15_tpGCLKBUF;
wire nx14650z1_SQMUX_BLSBR3_tpGCLKBUF;
wire nx14855z2;
wire nx15998z1;
wire nx15998z1_CAND2_TLSTR_11_tpGCLKBUF;
wire nx15998z1_CAND2_TLSTR_12_tpGCLKBUF;
wire nx15998z1_CAND2_TLSTR_13_tpGCLKBUF;
wire nx15998z1_CAND2_TLSTR_14_tpGCLKBUF;
wire nx15998z1_SQMUX_TLSTR2_tpGCLKBUF;
wire nx16644z1;
wire nx16644z2;
wire nx1674z1;
wire nx17641z1;
wire nx1800z1;
wire nx18281z3;
wire nx18527z1;
wire nx18527z8;
wire nx19381z1;
wire nx19726z1;
wire nx20469z1;
wire nx20521z1;
wire nx20942z2;
wire nx21518z1;
wire nx22012z2;
wire nx22245z1;
wire nx22245z2;
wire nx22245z2_CAND2_BLSBL_5_tpGCLKBUF;
wire nx22245z2_CAND2_BLSBL_6_tpGCLKBUF;
wire nx22245z2_CAND2_BLSBL_7_tpGCLKBUF;
wire nx22245z2_CAND2_BLSBL_8_tpGCLKBUF;
wire nx22245z2_CAND2_BLSTL_5_tpGCLKBUF;
wire nx22245z2_CAND2_BLSTL_6_tpGCLKBUF;
wire nx22245z2_CAND2_BLSTL_7_tpGCLKBUF;
wire nx22245z2_CAND2_BLSTL_8_tpGCLKBUF;
wire nx22245z2_QMUX_BL2_tpGCLKBUF;
wire nx22245z2_SQMUX_BLSBL2_tpGCLKBUF;
wire nx22245z2_SQMUX_BLSTL2_tpGCLKBUF;
wire nx22515z1;
wire nx23147z1;
wire nx25587z1;
wire nx25587z2;
wire nx25587z2_CAND2_TRSTR_25_tpGCLKBUF;
wire nx25587z2_CAND2_TRSTR_26_tpGCLKBUF;
wire nx25587z2_SQMUX_TRSTR2_tpGCLKBUF;
wire nx25788z3;
wire nx25788z3_CAND4_BRSBR_25_tpGCLKBUF;
wire nx25788z3_CAND4_BRSBR_26_tpGCLKBUF;
wire nx25788z3_CAND4_BRSBR_27_tpGCLKBUF;
wire nx25788z3_CAND4_BRSBR_28_tpGCLKBUF;
wire nx25788z3_CAND4_BRSBR_29_tpGCLKBUF;
wire nx25788z3_SQMUX_BRSBR4_tpGCLKBUF;
wire nx28356z1;
wire nx30664z1;
wire nx30923z2;
wire nx32122z1;
wire nx32231z2;
wire nx32231z2_CAND4_TLSTR_14_tpGCLKBUF;
wire nx32231z2_CAND4_TLSTR_15_tpGCLKBUF;
wire nx32231z2_SQMUX_TLSTR4_tpGCLKBUF;
wire nx33579z1;
wire nx33579z1_CAND2_BLSBR_11_tpGCLKBUF;
wire nx33579z1_CAND2_BLSBR_12_tpGCLKBUF;
wire nx33579z1_CAND2_BLSBR_13_tpGCLKBUF;
wire nx33579z1_CAND2_BLSBR_14_tpGCLKBUF;
wire nx33579z1_SQMUX_BLSBR2_tpGCLKBUF;
wire nx34006z1;
wire nx34006z2;
wire nx34006z2_CAND2_TLSTL_4_tpGCLKBUF;
wire nx34006z2_CAND2_TLSTL_5_tpGCLKBUF;
wire nx34006z2_CAND2_TLSTL_6_tpGCLKBUF;
wire nx34006z2_CAND2_TLSTL_7_tpGCLKBUF;
wire nx34006z2_CAND2_TLSTL_8_tpGCLKBUF;
wire nx34006z2_SQMUX_TLSTL2_tpGCLKBUF;
wire nx34850z5;
wire nx35588z2;
wire nx36058z2;
wire nx36058z2_CAND4_TRSTR_25_tpGCLKBUF;
wire nx36058z2_CAND4_TRSTR_26_tpGCLKBUF;
wire nx36058z2_CAND4_TRSTR_27_tpGCLKBUF;
wire nx36058z2_CAND4_TRSTR_28_tpGCLKBUF;
wire nx36058z2_CAND4_TRSTR_29_tpGCLKBUF;
wire nx36058z2_CAND5_TRSBR_25_tpGCLKBUF;
wire nx36058z2_CAND5_TRSBR_26_tpGCLKBUF;
wire nx36058z2_CAND5_TRSBR_27_tpGCLKBUF;
wire nx36058z2_CAND5_TRSBR_28_tpGCLKBUF;
wire nx36058z2_CAND5_TRSBR_29_tpGCLKBUF;
wire nx36058z2_SQMUX_TRSBR5_tpGCLKBUF;
wire nx36058z2_SQMUX_TRSTR4_tpGCLKBUF;
wire nx3668z1;
wire nx3668z8;
wire nx36808z2;
wire nx36875z1;
wire nx3786z2;
wire nx3786z2_CAND5_BRSBR_25_tpGCLKBUF;
wire nx3786z2_CAND5_BRSBR_26_tpGCLKBUF;
wire nx3786z2_CAND5_BRSBR_27_tpGCLKBUF;
wire nx3786z2_SQMUX_BRSBR5_tpGCLKBUF;
wire nx3850z2;
wire nx3850z2_CAND3_BRSBL_23_tpGCLKBUF;
wire nx3850z2_CAND3_BRSBL_24_tpGCLKBUF;
wire nx3850z2_CAND3_BRSBR_25_tpGCLKBUF;
wire nx3850z2_CAND3_BRSBR_26_tpGCLKBUF;
wire nx3850z2_CAND3_BRSBR_27_tpGCLKBUF;
wire nx3850z2_QMUX_BR3_tpGCLKBUF;
wire nx3850z2_SQMUX_BRSBL3_tpGCLKBUF;
wire nx3850z2_SQMUX_BRSBR3_tpGCLKBUF;
wire nx39177z2;
wire nx39177z2_CAND5_TRSTR_25_tpGCLKBUF;
wire nx39177z2_CAND5_TRSTR_26_tpGCLKBUF;
wire nx39177z2_SQMUX_TRSTR5_tpGCLKBUF;
wire nx39673z1;
wire nx39673z6;
wire nx39840z1;
wire nx39840z1_CAND4_TLSTL_1_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_2_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_3_tpGCLKBUF;
wire nx39840z1_CAND4_TLSTL_4_tpGCLKBUF;
wire nx39840z1_SQMUX_TLSTL4_tpGCLKBUF;
wire nx40545z1;
wire nx40546z1;
wire nx40547z1;
wire nx40548z1;
wire nx40548z2;
wire nx40548z2_CAND3_BRSTR_25_tpGCLKBUF;
wire nx40548z2_CAND3_BRSTR_26_tpGCLKBUF;
wire nx40548z2_CAND3_BRSTR_27_tpGCLKBUF;
wire nx40548z2_SQMUX_BRSTR3_tpGCLKBUF;
wire nx40728z1;
wire nx41096z1;
wire nx41097z1;
wire nx41193z2;
wire nx41193z2_CAND3_TRSTL_17_tpGCLKBUF;
wire nx41193z2_CAND3_TRSTL_18_tpGCLKBUF;
wire nx41193z2_CAND3_TRSTL_19_tpGCLKBUF;
wire nx41193z2_CAND3_TRSTL_20_tpGCLKBUF;
wire nx41193z2_CAND3_TRSTL_21_tpGCLKBUF;
wire nx41193z2_SQMUX_TRSTL3_tpGCLKBUF;
wire nx41667z1;
wire nx42281z2;
wire nx42664z1;
wire nx42928z2;
wire nx42928z2_CAND3_TLSTL_4_tpGCLKBUF;
wire nx42928z2_CAND3_TLSTL_5_tpGCLKBUF;
wire nx42928z2_CAND3_TLSTL_6_tpGCLKBUF;
wire nx42928z2_CAND3_TLSTL_7_tpGCLKBUF;
wire nx42928z2_CAND3_TLSTL_8_tpGCLKBUF;
wire nx42928z2_SQMUX_TLSTL3_tpGCLKBUF;
wire nx43661z1;
wire nx44608z1;
wire nx44608z1_CAND2_TLSBL_1_tpGCLKBUF;
wire nx44608z1_CAND2_TLSBL_2_tpGCLKBUF;
wire nx44608z1_CAND2_TLSBL_3_tpGCLKBUF;
wire nx44608z1_CAND2_TLSBL_4_tpGCLKBUF;
wire nx44608z1_CAND2_TLSBL_5_tpGCLKBUF;
wire nx44608z1_SQMUX_TLSBL2_tpGCLKBUF;
wire nx45272z2;
wire nx46309z2;
wire nx48658z2;
wire nx4939z1;
wire nx4939z1_CAND3_BLSTL_1_tpGCLKBUF;
wire nx4939z1_CAND3_BLSTL_2_tpGCLKBUF;
wire nx4939z1_CAND3_BLSTL_3_tpGCLKBUF;
wire nx4939z1_CAND3_BLSTL_4_tpGCLKBUF;
wire nx4939z1_CAND3_BLSTL_5_tpGCLKBUF;
wire nx4939z1_SQMUX_BLSTL3_tpGCLKBUF;
wire nx49703z1;
wire nx49808z66;
wire nx49871z1;
wire nx50994z1;
wire nx50994z2;
wire nx50995z1;
wire nx50995z3;
wire nx50996z1;
wire nx50996z2;
wire nx50997z1;
wire nx50997z2;
wire nx53524z1;
wire nx56739z2;
wire nx57183z1;
wire nx58292z1;
wire nx58361z1;
wire nx58678z1;
wire nx60509z1;
wire nx60851z2;
wire nx60851z2_CAND4_BRSTR_27_tpGCLKBUF;
wire nx60851z2_CAND4_BRSTR_28_tpGCLKBUF;
wire nx60851z2_SQMUX_BRSTR4_tpGCLKBUF;
wire nx60936z2;
wire nx60936z2_CAND5_BRSTR_25_tpGCLKBUF;
wire nx60936z2_CAND5_BRSTR_26_tpGCLKBUF;
wire nx60936z2_CAND5_BRSTR_27_tpGCLKBUF;
wire nx60936z2_SQMUX_BRSTR5_tpGCLKBUF;
wire nx63842z2;
wire nx63842z2_CAND1_BRSTR_25_tpGCLKBUF;
wire nx63842z2_CAND1_BRSTR_26_tpGCLKBUF;
wire nx63842z2_CAND1_BRSTR_27_tpGCLKBUF;
wire nx63842z2_CAND1_BRSTR_28_tpGCLKBUF;
wire nx63842z2_SQMUX_BRSTR1_tpGCLKBUF;
wire nx64401z2;
wire nx65216z1;
wire nx677z1;
wire nx7012z1;
wire nx7012z2;
wire nx9707z1;
wire nx9707z1_CAND5_BLSTL_1_tpGCLKBUF;
wire nx9707z1_CAND5_BLSTL_2_tpGCLKBUF;
wire nx9707z1_CAND5_BLSTL_3_tpGCLKBUF;
wire nx9707z1_CAND5_BLSTL_5_tpGCLKBUF;
wire nx9707z1_SQMUX_BLSTL5_tpGCLKBUF;
wire p0_fsm_0__CAND5_TLSTL_7_tpGCLKBUF;
wire p0_fsm_0__CAND5_TLSTL_8_tpGCLKBUF;
wire p0_fsm_0__SQMUX_TLSTL5_tpGCLKBUF;
wire p1_fsm_0__CAND4_TRSTL_22_tpGCLKBUF;
wire p1_fsm_0__CAND4_TRSTL_23_tpGCLKBUF;
wire p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF;
wire p1_fsm_0__SQMUX_TRSTL4_tpGCLKBUF;
wire p2_fsm_0__CAND4_BLSBL_6_tpGCLKBUF;
wire p2_fsm_0__CAND4_BLSBL_7_tpGCLKBUF;
wire p2_fsm_0__CAND4_BLSBL_8_tpGCLKBUF;
wire p2_fsm_0__SQMUX_BLSBL4_tpGCLKBUF;
wire p2_fsm_4__CAND5_BLSBL_5_tpGCLKBUF;
wire p2_fsm_4__CAND5_BLSBL_6_tpGCLKBUF;
wire p2_fsm_4__CAND5_BLSBL_8_tpGCLKBUF;
wire p2_fsm_4__SQMUX_BLSBL5_tpGCLKBUF;
wire p3_fsm_0__CAND1_BRSBL_21_tpGCLKBUF;
wire p3_fsm_0__CAND1_BRSBL_22_tpGCLKBUF;
wire p3_fsm_0__CAND1_BRSBL_23_tpGCLKBUF;
wire p3_fsm_0__CAND1_BRSBL_24_tpGCLKBUF;
wire p3_fsm_0__SQMUX_BRSBL1_tpGCLKBUF;
wire saved_REQ;
wire tcdm_clk_p0;
wire tcdm_clk_p1;
wire tcdm_clk_p2;
wire tcdm_clk_p3;
wire tcdm_fmo_p0;
wire tcdm_fmo_p0_int;
wire tcdm_fmo_p1;
wire tcdm_fmo_p1_int;
wire tcdm_fmo_p2;
wire tcdm_fmo_p2_int;
wire tcdm_fmo_p3;
wire tcdm_fmo_p3_int;
wire tcdm_gnt_p0;
wire tcdm_gnt_p0_int;
wire tcdm_gnt_p1;
wire tcdm_gnt_p1_int;
wire tcdm_gnt_p2;
wire tcdm_gnt_p2_int;
wire tcdm_gnt_p3;
wire tcdm_gnt_p3_int;
wire tcdm_req_p0;
wire tcdm_req_p0_dup_0;
wire tcdm_req_p1;
wire tcdm_req_p1_dup_0;
wire tcdm_req_p2;
wire tcdm_req_p2_dup_0;
wire tcdm_req_p3;
wire tcdm_req_p3_dup_0;
wire tcdm_valid_p0;
wire tcdm_valid_p0_int;
wire tcdm_valid_p0_int_CAND3_TLSTR_10_tpGCLKBUF;
wire tcdm_valid_p0_int_CAND3_TLSTR_13_tpGCLKBUF;
wire tcdm_valid_p0_int_CAND3_TLSTR_14_tpGCLKBUF;
wire tcdm_valid_p0_int_CAND3_TLSTR_15_tpGCLKBUF;
wire tcdm_valid_p0_int_CAND3_TLSTR_16_tpGCLKBUF;
wire tcdm_valid_p0_int_CAND3_TLSTR_9_tpGCLKBUF;
wire tcdm_valid_p0_int_SQMUX_TLSTR3_tpGCLKBUF;
wire tcdm_valid_p1;
wire tcdm_valid_p1_int;
wire tcdm_valid_p2;
wire tcdm_valid_p2_int;
wire tcdm_valid_p2_int_CAND2_BLSTR_10_tpGCLKBUF;
wire tcdm_valid_p2_int_CAND2_BLSTR_12_tpGCLKBUF;
wire tcdm_valid_p2_int_CAND2_BLSTR_13_tpGCLKBUF;
wire tcdm_valid_p2_int_CAND2_BLSTR_15_tpGCLKBUF;
wire tcdm_valid_p2_int_SQMUX_BLSTR2_tpGCLKBUF;
wire tcdm_valid_p3;
wire tcdm_valid_p3_int;
wire tcdm_wen_p0;
wire tcdm_wen_p0_dup_0;
wire tcdm_wen_p1;
wire tcdm_wen_p1_dup_0;
wire tcdm_wen_p2;
wire tcdm_wen_p2_dup_0;
wire tcdm_wen_p3;
wire tcdm_wen_p3_dup_0;
wire [5:0] CLK;
wire [5:0] CLK_int;
wire [3:0] RESET;
wire [3:0] RESET_int;
wire [1:0] apb_fsm;
wire [2:0] cnt1;
wire [2:0] cnt2;
wire [2:0] cnt3;
wire [2:0] cnt4;
wire [2:0] cnt5;
wire [31:0] control_in;
wire [31:0] control_in_int;
wire [15:0] events_o;
wire [79:0] fpgaio_in;
wire [79:0] fpgaio_in_int;
wire [79:0] fpgaio_oe;
wire [79:0] fpgaio_oe_dup_0;
wire [79:0] fpgaio_out;
wire [79:0] fpgaio_out_dup_0;
wire [15:0] i_events;
wire [3:0] last_control;
wire [19:0] lint_ADDR;
wire [19:0] lint_ADDR_int;
wire [3:0] lint_BE;
wire [3:0] lint_BE_int;
wire [31:0] lint_RDATA;
wire [31:0] lint_RDATA_dup_0;
wire [31:0] lint_WDATA;
wire [31:0] lint_WDATA_int;
wire [11:0] m0_coef_raddr;
wire [11:0] m0_coef_raddr_dup_0;
wire [31:0] m0_coef_rdata;
wire [31:0] m0_coef_rdata_int;
wire [1:0] m0_coef_rmode;
wire [1:0] m0_coef_rmode_dup_0;
wire [11:0] m0_coef_waddr;
wire [11:0] m0_coef_waddr_dup_0;
wire [31:0] m0_coef_wdata;
wire [31:0] m0_coef_wdata_dup_0;
wire [1:0] m0_coef_wmode;
wire [1:0] m0_coef_wmode_dup_0;
wire [31:0] m0_m0_coef_in;
wire [30:7] m0_m0_control;
wire [31:0] m0_m0_dataout;
wire [31:0] m0_m0_dataout_int;
wire [1:0] m0_m0_mode;
wire [1:0] m0_m0_mode_dup_0;
wire [31:0] m0_m0_oper_in;
wire [5:0] m0_m0_outsel;
wire [5:0] m0_m0_outsel_dup_0;
wire [31:0] m0_m1_coef_in;
wire [30:7] m0_m1_control;
wire [31:0] m0_m1_dataout;
wire [31:0] m0_m1_dataout_int;
wire [1:0] m0_m1_mode;
wire [1:0] m0_m1_mode_dup_0;
wire [31:0] m0_m1_oper_in;
wire [5:0] m0_m1_outsel;
wire [5:0] m0_m1_outsel_dup_0;
wire [11:0] m0_oper0_raddr;
wire [11:0] m0_oper0_raddr_dup_0;
wire [31:0] m0_oper0_rdata;
wire [31:0] m0_oper0_rdata_int;
wire [1:0] m0_oper0_rmode;
wire [1:0] m0_oper0_rmode_dup_0;
wire [11:0] m0_oper0_waddr;
wire [11:0] m0_oper0_waddr_dup_0;
wire [31:0] m0_oper0_wdata;
wire [31:0] m0_oper0_wdata_dup_0;
wire [1:0] m0_oper0_wmode;
wire [1:0] m0_oper0_wmode_dup_0;
wire [11:0] m0_oper1_raddr;
wire [11:0] m0_oper1_raddr_dup_0;
wire [31:0] m0_oper1_rdata;
wire [31:0] m0_oper1_rdata_int;
wire [1:0] m0_oper1_rmode;
wire [1:0] m0_oper1_rmode_dup_0;
wire [11:0] m0_oper1_waddr;
wire [11:0] m0_oper1_waddr_dup_0;
wire [31:0] m0_oper1_wdata;
wire [31:0] m0_oper1_wdata_dup_0;
wire [1:0] m0_oper1_wmode;
wire [1:0] m0_oper1_wmode_dup_0;
wire [31:15] m0_ram_control;
wire [11:0] m1_coef_raddr;
wire [11:0] m1_coef_raddr_dup_0;
wire [31:0] m1_coef_rdata;
wire [31:0] m1_coef_rdata_int;
wire [1:0] m1_coef_rmode;
wire [1:0] m1_coef_rmode_dup_0;
wire [11:0] m1_coef_waddr;
wire [11:0] m1_coef_waddr_dup_0;
wire [31:0] m1_coef_wdata;
wire [31:0] m1_coef_wdata_dup_0;
wire [1:0] m1_coef_wmode;
wire [1:0] m1_coef_wmode_dup_0;
wire [31:0] m1_m0_coef_in;
wire [30:7] m1_m0_control;
wire [31:0] m1_m0_dataout;
wire [31:0] m1_m0_dataout_int;
wire [1:0] m1_m0_mode;
wire [1:0] m1_m0_mode_dup_0;
wire [31:0] m1_m0_oper_in;
wire [5:0] m1_m0_outsel;
wire [5:0] m1_m0_outsel_dup_0;
wire [31:0] m1_m1_coef_in;
wire [30:0] m1_m1_control;
wire [31:0] m1_m1_dataout;
wire [31:0] m1_m1_dataout_int;
wire [1:0] m1_m1_mode;
wire [1:0] m1_m1_mode_dup_0;
wire [31:0] m1_m1_oper_in;
wire [5:0] m1_m1_outsel;
wire [11:0] m1_oper0_raddr;
wire [11:2] m1_oper0_raddr_dup_0;
wire [31:0] m1_oper0_rdata;
wire [31:0] m1_oper0_rdata_int;
wire [1:0] m1_oper0_rmode;
wire [1:0] m1_oper0_rmode_dup_0;
wire [11:0] m1_oper0_waddr;
wire [11:0] m1_oper0_waddr_dup_0;
wire [31:0] m1_oper0_wdata;
wire [31:0] m1_oper0_wdata_dup_0;
wire [1:0] m1_oper0_wmode;
wire [1:0] m1_oper0_wmode_dup_0;
wire [11:0] m1_oper1_raddr;
wire [11:2] m1_oper1_raddr_dup_0;
wire [31:0] m1_oper1_rdata;
wire [31:0] m1_oper1_rdata_int;
wire [1:0] m1_oper1_rmode;
wire [1:0] m1_oper1_rmode_dup_0;
wire [11:0] m1_oper1_waddr;
wire [11:0] m1_oper1_waddr_dup_0;
wire [31:0] m1_oper1_wdata;
wire [31:0] m1_oper1_wdata_dup_0;
wire [1:0] m1_oper1_wmode;
wire [1:0] m1_oper1_wmode_dup_0;
wire [31:15] m1_ram_control;
wire [11:0] p0_cnt;
wire [4:0] p0_fsm;
wire [11:0] p1_cnt;
wire [4:0] p1_fsm;
wire [11:0] p2_cnt;
wire [4:0] p2_fsm;
wire [11:0] p3_cnt;
wire [4:0] p3_fsm;
wire [31:0] status_out;
wire [19:0] tcdm_addr_p0;
wire [19:0] tcdm_addr_p0_dup_0;
wire [19:0] tcdm_addr_p1;
wire [19:0] tcdm_addr_p1_dup_0;
wire [19:0] tcdm_addr_p2;
wire [19:0] tcdm_addr_p2_dup_0;
wire [19:0] tcdm_addr_p3;
wire [19:0] tcdm_addr_p3_dup_0;
wire [3:0] tcdm_be_p0;
wire [3:0] tcdm_be_p0_17n77s1;
wire [3:0] tcdm_be_p0_dup_0;
wire [3:0] tcdm_be_p1;
wire [3:0] tcdm_be_p1_dup_0;
wire [3:0] tcdm_be_p2;
wire [3:0] tcdm_be_p2_dup_0;
wire [3:0] tcdm_be_p3;
wire [3:0] tcdm_be_p3_dup_0;
wire [31:0] tcdm_rdata_p0;
wire [31:0] tcdm_rdata_p0_int;
wire [31:0] tcdm_rdata_p1;
wire [31:0] tcdm_rdata_p1_int;
wire [31:0] tcdm_rdata_p2;
wire [31:0] tcdm_rdata_p2_int;
wire [31:0] tcdm_rdata_p3;
wire [31:0] tcdm_rdata_p3_int;
wire [31:0] tcdm_result_p0;
wire [31:0] tcdm_result_p1;
wire [31:0] tcdm_result_p2;
wire [31:0] tcdm_result_p3;
wire [31:0] tcdm_wdata_p0;
wire [31:0] tcdm_wdata_p0_dup_0;
wire [31:0] tcdm_wdata_p1;
wire [31:0] tcdm_wdata_p1_dup_0;
wire [31:0] tcdm_wdata_p2;
wire [31:0] tcdm_wdata_p2_dup_0;
wire [31:0] tcdm_wdata_p3;
wire [31:0] tcdm_wdata_p3_dup_0;
wire [7:0] version;

	LOGIC_0 QL_INST_A6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx39840z1_CAND4_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx39840z1_CAND4_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx39840z1_CAND4_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx39840z1_CAND4_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx39840z1_CAND4_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[26]),.Q1EN(nx39840z1_CAND4_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx39840z1_CAND4_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx39840z1_CAND4_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A8_0 (.tFragBitInfo(16'b1111011111110111),.bFragBitInfo(16'b1111000011110111),.B0I0(fpgaio_oe_dup_0[22]),.B0I1(NET_75),.B0I2(lint_ADDR_int[11]),.B0I3(NET_73),.CD0S(VCC),.Q0DI(lint_WDATA_int[22]),.Q0EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_oe_dup_0[22]),.T0I1(NET_75),.T0I2(lint_ADDR_int[11]),.T0I3(NET_73),.TB0S(fpgaio_out_dup_0[22]),.C0Z(NET_554),.Q0Z(fpgaio_oe_dup_0[22]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A8_1 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.T1I0(NET_73),.T1I1(fpgaio_out_dup_0[7]),.T1I2(lint_ADDR_int[11]),.T1I3(GND),.C1Z(NET_607),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_A8_2 (.tFragBitInfo(16'b1111001111111111),.bFragBitInfo(16'b1111000111110101),.B2I0(fpgaio_out_dup_0[21]),.B2I1(NET_75),.B2I2(lint_ADDR_int[11]),.B2I3(fpgaio_oe_dup_0[21]),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_out_dup_0[21]),.T2I1(NET_75),.T2I2(lint_ADDR_int[11]),.T2I3(fpgaio_oe_dup_0[21]),.TB2S(NET_73),.C2Z(NET_922),.Q2Z(fpgaio_oe_dup_0[21]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_A8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx39840z1_CAND4_TLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_1_padClk),.QRT(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A9_0 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int_11__CAND4_TLSBL_1_tpGCLKBUF),.T0I1(fpgaio_out_dup_0[12]),.T0I2(GND),.T0I3(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.TB0S(GND),.C0Z(NET_321),.Q0Z(fpgaio_oe_dup_0[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[13]),.Q2EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A9_3 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int_11__CAND4_TLSBL_1_tpGCLKBUF),.T3I1(GND),.T3I2(fpgaio_out_dup_0[26]),.T3I3(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.TB3S(GND),.C3Z(NET_657),.Q3Z(fpgaio_out_dup_0[31]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_A10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001000),.B0I0(fpgaio_out_dup_0[0]),.B0I1(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.B0I2(GND),.B0I3(lint_ADDR_int_11__CAND4_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.B0Z(NET_132),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000001000000),.B2I0(GND),.B2I1(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.B2I2(fpgaio_out_dup_0[17]),.B2I3(lint_ADDR_int_11__CAND4_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.B2Z(NET_447),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A13_0 (.tFragBitInfo(16'b0000011100000111),.bFragBitInfo(16'b0000000000000111),.B0I0(NET_133),.B0I1(fpgaio_out_dup_0[39]),.B0I2(NET_607),.B0I3(fpgaio_oe_dup_0[7]),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(NET_133),.T0I1(fpgaio_out_dup_0[39]),.T0I2(NET_607),.T0I3(fpgaio_oe_dup_0[7]),.TB0S(NET_134),.C0Z(NET_590),.Q0Z(fpgaio_oe_dup_0[7]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A13_1 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int_11__CAND4_TLSBL_1_tpGCLKBUF),.T1I1(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.T1I2(GND),.T1I3(fpgaio_out_dup_0[2]),.C1Z(NET_909),.Q1Z(fpgaio_oe_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_A13_2 (.tFragBitInfo(16'b0001000100110011),.bFragBitInfo(16'b0000000100000011),.B2I0(NET_133),.B2I1(NET_132),.B2I2(fpgaio_oe_dup_0[0]),.B2I3(fpgaio_out_dup_0[32]),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T2I0(NET_133),.T2I1(NET_132),.T2I2(fpgaio_oe_dup_0[0]),.T2I3(fpgaio_out_dup_0[32]),.TB2S(NET_134),.C2Z(NET_94),.Q2Z(fpgaio_oe_dup_0[9]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_A13_3 (.tFragBitInfo(16'b0001001100010011),.bFragBitInfo(16'b0000000000010011),.B3I0(NET_133),.B3I1(fpgaio_oe_dup_0[2]),.B3I2(fpgaio_out_dup_0[34]),.B3I3(NET_909),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_out_dup_0[34]),.T3I1(NET_909),.T3I2(NET_133),.T3I3(fpgaio_oe_dup_0[2]),.TB3S(NET_134),.C3Z(NET_892),.Q3Z(fpgaio_oe_dup_0[4]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_A14_0 (.tFragBitInfo(16'b0000010100001111),.bFragBitInfo(16'b0000000100000011),.B0I0(fpgaio_oe_dup_0[58]),.B0I1(fpgaio_oe_dup_0[26]),.B0I2(NET_657),.B0I3(NET_146),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_oe_dup_0[58]),.T0I1(fpgaio_oe_dup_0[26]),.T0I2(NET_657),.T0I3(NET_146),.TB0S(NET_134),.C0Z(NET_654),.Q0Z(fpgaio_oe_dup_0[13]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A14_1 (.tFragBitInfo(16'b0000011100000111),.bFragBitInfo(16'b0000000100010001),.B1I0(NET_321),.B1I1(fpgaio_oe_dup_0[12]),.B1I2(fpgaio_out_dup_0[44]),.B1I3(NET_133),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[44]),.T1I1(NET_133),.T1I2(NET_321),.T1I3(fpgaio_oe_dup_0[12]),.TB1S(NET_134),.C1Z(NET_304),.Q1Z(fpgaio_oe_dup_0[10]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_A14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000010000000000),.B2I0(GND),.B2I1(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.B2I2(lint_ADDR_int_11__CAND4_TLSBL_1_tpGCLKBUF),.B2I3(fpgaio_out_dup_0[29]),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.B2Z(NET_722),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A14_3 (.tFragBitInfo(16'b0001000101010101),.bFragBitInfo(16'b0000000100000101),.B3I0(fpgaio_oe_dup_0[29]),.B3I1(fpgaio_oe_dup_0[61]),.B3I2(NET_722),.B3I3(NET_146),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T3I0(NET_722),.T3I1(NET_146),.T3I2(fpgaio_oe_dup_0[29]),.T3I3(fpgaio_oe_dup_0[61]),.TB3S(NET_134),.C3Z(NET_719),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_A15_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.B0I1(NET_72),.B0I2(fpgaio_out_dup_0[31]),.B0I3(fpgaio_oe_dup_0[63]),.T0I0(fpgaio_out_dup_0[40]),.T0I1(fpgaio_oe_dup_0[8]),.T0I2(NET_76),.T0I3(NET_75_CAND5_TLSBL_1_tpGCLKBUF),.TB0S(GND),.B0Z(NET_772),.C0Z(NET_384),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_A15_1 (.tFragBitInfo(16'b0000110011001100),.bFragBitInfo(16'b0000011100000000),.B1I0(fpgaio_oe_dup_0[31]),.B1I1(NET_75_CAND5_TLSBL_1_tpGCLKBUF),.B1I2(fpgaio_out_dup_0[63]),.B1I3(NET_772),.T1I0(fpgaio_out_dup_0[63]),.T1I1(NET_772),.T1I2(fpgaio_oe_dup_0[31]),.T1I3(NET_75_CAND5_TLSBL_1_tpGCLKBUF),.TB1S(NET_76),.C1Z(NET_773),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_A15_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.B2I1(fpgaio_out_dup_0[20]),.B2I2(NET_76),.B2I3(fpgaio_out_dup_0[52]),.T2I0(lint_ADDR_int[16]),.T2I1(lint_ADDR_int[18]),.T2I2(lint_ADDR_int[19]),.T2I3(lint_ADDR_int[17]),.TB2S(GND),.B2Z(NET_520),.C2Z(NET_9),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_A15_3 (.tFragBitInfo(16'b0010001010101010),.bFragBitInfo(16'b0001000001010000),.B3I0(fpgaio_out_dup_0[8]),.B3I1(fpgaio_oe_dup_0[40]),.B3I2(NET_384),.B3I3(NET_72),.T3I0(NET_384),.T3I1(NET_72),.T3I2(fpgaio_out_dup_0[8]),.T3I3(fpgaio_oe_dup_0[40]),.TB3S(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.C3Z(NET_376),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_A16_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_oe_dup_0[4]),.B0I1(fpgaio_out_dup_0[36]),.B0I2(NET_75_CAND5_TLSBL_1_tpGCLKBUF),.B0I3(NET_76),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T0I0(NET_76),.T0I1(fpgaio_out_dup_0[45]),.T0I2(NET_75_CAND5_TLSBL_1_tpGCLKBUF),.T0I3(fpgaio_oe_dup_0[13]),.TB0S(GND),.B0Z(NET_856),.C0Z(NET_338),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A16_1 (.tFragBitInfo(16'b0100010011001100),.bFragBitInfo(16'b0001010100000000),.B1I0(fpgaio_out_dup_0[4]),.B1I1(fpgaio_oe_dup_0[36]),.B1I2(NET_72),.B1I3(NET_856),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T1I0(NET_72),.T1I1(NET_856),.T1I2(fpgaio_out_dup_0[4]),.T1I3(fpgaio_oe_dup_0[36]),.TB1S(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.C1Z(NET_857),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_A16_2 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0000000000101010),.B2I0(NET_338),.B2I1(NET_72),.B2I2(fpgaio_oe_dup_0[45]),.B2I3(fpgaio_out_dup_0[13]),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx9707z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.T2I0(NET_338),.T2I1(NET_72),.T2I2(fpgaio_oe_dup_0[45]),.T2I3(fpgaio_out_dup_0[13]),.TB2S(NET_73_CAND3_TLSBL_1_tpGCLKBUF),.C2Z(NET_339),.Q2Z(fpgaio_oe_dup_0[37]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_A16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx9707z1),.QCK(CLK_int_0__CAND0_TLSBL_1_padClk),.QRT(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[58]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A17_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_75),.B0I1(NET_76),.B0I2(fpgaio_out_dup_0[42]),.B0I3(fpgaio_oe_dup_0[10]),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T0I0(NET_75),.T0I1(NET_76),.T0I2(fpgaio_oe_dup_0[9]),.T0I3(fpgaio_out_dup_0[41]),.TB0S(GND),.B0Z(NET_269),.C0Z(NET_239),.Q0Z(fpgaio_oe_dup_0[56]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A17_1 (.tFragBitInfo(16'b0101111100000000),.bFragBitInfo(16'b0000000001001100),.B1I0(NET_72),.B1I1(NET_269),.B1I2(fpgaio_oe_dup_0[42]),.B1I3(fpgaio_out_dup_0[10]),.CD1S(VCC),.Q1DI(lint_WDATA_int[4]),.Q1EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_oe_dup_0[42]),.T1I1(fpgaio_out_dup_0[10]),.T1I2(NET_72),.T1I3(NET_269),.TB1S(NET_73),.C1Z(NET_261),.Q1Z(fpgaio_oe_dup_0[36]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_A17_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_75),.B2I1(NET_72),.B2I2(fpgaio_oe_dup_0[57]),.B2I3(fpgaio_oe_dup_0[25]),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(NET_73),.T2I1(fpgaio_out_dup_0[11]),.T2I2(fpgaio_out_dup_0[43]),.T2I3(NET_76),.TB2S(GND),.B2Z(NET_642),.C2Z(NET_285),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_A17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[45]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[63]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[49]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A18_2 (.tFragBitInfo(16'b0001010100010101),.bFragBitInfo(16'b0000000000010101),.B2I0(NET_447),.B2I1(NET_146),.B2I2(fpgaio_oe_dup_0[49]),.B2I3(fpgaio_out_dup_0[49]),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(NET_447),.T2I1(NET_146),.T2I2(fpgaio_oe_dup_0[49]),.T2I3(fpgaio_out_dup_0[49]),.TB2S(NET_133),.C2Z(NET_438),.Q2Z(fpgaio_oe_dup_0[61]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_A18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[35]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[40]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[63]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[34]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[42]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A20_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_oe_dup_0[53]),.T0I1(NET_146),.T0I2(NET_133),.T0I3(fpgaio_out_dup_0[53]),.TB0S(GND),.C0Z(NET_531),.Q0Z(fpgaio_oe_dup_0[57]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_A20_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T1I0(NET_146),.T1I1(fpgaio_out_dup_0[54]),.T1I2(NET_133),.T1I3(fpgaio_oe_dup_0[54]),.TB1S(GND),.C1Z(NET_555),.Q1Z(fpgaio_oe_dup_0[54]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_A20_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_146),.B2I1(fpgaio_out_dup_0[55]),.B2I2(NET_133),.B2I3(fpgaio_oe_dup_0[55]),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_oe_dup_0[50]),.T2I1(NET_146),.T2I2(NET_133),.T2I3(fpgaio_out_dup_0[50]),.TB2S(GND),.B2Z(NET_573),.C2Z(NET_460),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_A20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[40]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[44]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[49]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[43]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[50]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[44]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[23]),.Q1EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[55]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[53]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[41]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[50]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[21]),.Q1EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[53]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[36]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[45]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[42]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[54]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[39]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_1_padClk),.QRT(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[57]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_A25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[55]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_A25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[52]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_A25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_A25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_1_padClk),.QRT(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx39840z1_CAND4_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx39840z1_CAND4_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx39840z1_CAND4_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx39840z1_CAND4_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[25]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx39840z1_CAND4_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx39840z1_CAND4_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B8_1 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(lint_ADDR_int[11]),.T1I2(NET_73),.T1I3(fpgaio_out_dup_0[6]),.C1Z(NET_807),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_B8_2 (.tFragBitInfo(16'b1111111101011111),.bFragBitInfo(16'b1111111100010011),.B2I0(NET_75),.B2I1(fpgaio_out_dup_0[23]),.B2I2(fpgaio_oe_dup_0[23]),.B2I3(lint_ADDR_int[11]),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx39840z1_CAND4_TLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.T2I0(NET_75),.T2I1(fpgaio_out_dup_0[23]),.T2I2(fpgaio_oe_dup_0[23]),.T2I3(lint_ADDR_int[11]),.TB2S(NET_73),.C2Z(NET_923),.Q2Z(fpgaio_out_dup_0[24]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_B8_3 (.tFragBitInfo(16'b1101110111111111),.bFragBitInfo(16'b1111111100010101),.B3I0(fpgaio_out_dup_0[18]),.B3I1(fpgaio_oe_dup_0[18]),.B3I2(NET_75),.B3I3(lint_ADDR_int[11]),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSTL_2_padClk),.QRT(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF),.QST(GND),.T3I0(NET_75),.T3I1(lint_ADDR_int[11]),.T3I2(fpgaio_out_dup_0[18]),.T3I3(fpgaio_oe_dup_0[18]),.TB3S(NET_73),.C3Z(NET_919),.Q3Z(fpgaio_oe_dup_0[23]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_B9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[6]),.Q0EN(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[16]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B0I0(fpgaio_out_dup_0[24]),.B0I1(lint_ADDR_int_11__CAND4_TLSBL_2_tpGCLKBUF),.B0I2(GND),.B0I3(NET_73_CAND3_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.B0Z(NET_618),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B10_3 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_out_dup_0[28]),.T3I1(lint_ADDR_int_11__CAND4_TLSBL_2_tpGCLKBUF),.T3I2(GND),.T3I3(NET_73_CAND3_TLSBL_2_tpGCLKBUF),.C3Z(NET_699),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_B11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[19]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B11_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[19]),.T1I1(lint_ADDR_int_11__CAND4_TLSBL_2_tpGCLKBUF),.T1I2(NET_73_CAND3_TLSBL_2_tpGCLKBUF),.T1I3(GND),.C1Z(NET_495),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_B11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[28]),.Q0EN(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[28]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[5]),.Q0EN(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B13_1 (.tFragBitInfo(16'b0000001100001111),.bFragBitInfo(16'b0000000100000101),.B1I0(NET_807),.B1I1(NET_133),.B1I2(fpgaio_oe_dup_0[6]),.B1I3(fpgaio_out_dup_0[38]),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_oe_dup_0[6]),.T1I1(fpgaio_out_dup_0[38]),.T1I2(NET_807),.T1I3(NET_133),.TB1S(NET_134),.C1Z(NET_790),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_B13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B14_0 (.tFragBitInfo(16'b0001001100010011),.bFragBitInfo(16'b0000000000010011),.B0I0(fpgaio_oe_dup_0[56]),.B0I1(NET_618),.B0I2(NET_146),.B0I3(fpgaio_oe_dup_0[24]),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_oe_dup_0[56]),.T0I1(NET_618),.T0I2(NET_146),.T0I3(fpgaio_oe_dup_0[24]),.TB0S(NET_134),.C0Z(NET_615),.Q0Z(fpgaio_oe_dup_0[30]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_B14_1 (.tFragBitInfo(16'b0000000000111111),.bFragBitInfo(16'b0000000100000011),.B1I0(fpgaio_oe_dup_0[60]),.B1I1(NET_699),.B1I2(fpgaio_oe_dup_0[28]),.B1I3(NET_146),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_oe_dup_0[28]),.T1I1(NET_146),.T1I2(fpgaio_oe_dup_0[60]),.T1I3(NET_699),.TB1S(NET_134),.C1Z(NET_696),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_B14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000100),.B2I0(GND),.B2I1(NET_75_CAND5_TLSBL_2_tpGCLKBUF),.B2I2(GND),.B2I3(lint_ADDR_int_11__CAND4_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.B2Z(NET_134),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B15_0 (.tFragBitInfo(16'b0011000011110000),.bFragBitInfo(16'b0001000001010000),.B0I0(fpgaio_out_dup_0[3]),.B0I1(fpgaio_out_dup_0[35]),.B0I2(NET_879),.B0I3(NET_76),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.T0I0(fpgaio_out_dup_0[3]),.T0I1(fpgaio_out_dup_0[35]),.T0I2(NET_879),.T0I3(NET_76),.TB0S(NET_73_CAND3_TLSBL_2_tpGCLKBUF),.C0Z(NET_871),.Q0Z(fpgaio_oe_dup_0[16]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_B15_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.T1I0(NET_76),.T1I1(fpgaio_out_dup_0[47]),.T1I2(fpgaio_oe_dup_0[15]),.T1I3(NET_75_CAND5_TLSBL_2_tpGCLKBUF),.TB1S(GND),.C1Z(NET_405),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_B15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(fpgaio_oe_dup_0[35]),.B2I1(fpgaio_oe_dup_0[3]),.B2I2(NET_72),.B2I3(NET_75_CAND5_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.B2Z(NET_879),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B15_3 (.tFragBitInfo(16'b0011000011110000),.bFragBitInfo(16'b0000001000001010),.B3I0(NET_405),.B3I1(NET_72),.B3I2(fpgaio_out_dup_0[15]),.B3I3(fpgaio_oe_dup_0[47]),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_2_padClk),.QRT(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_out_dup_0[15]),.T3I1(fpgaio_oe_dup_0[47]),.T3I2(NET_405),.T3I3(NET_72),.TB3S(NET_73_CAND3_TLSBL_2_tpGCLKBUF),.C3Z(NET_397),.Q3Z(fpgaio_oe_dup_0[15]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_B16_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_73_CAND3_TLSBL_2_tpGCLKBUF),.B0I1(NET_72),.B0I2(fpgaio_out_dup_0[5]),.B0I3(fpgaio_oe_dup_0[37]),.T0I0(NET_73_CAND3_TLSBL_2_tpGCLKBUF),.T0I1(NET_72),.T0I2(fpgaio_out_dup_0[1]),.T0I3(fpgaio_oe_dup_0[33]),.TB0S(GND),.B0Z(NET_826),.C0Z(NET_11),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_B16_1 (.tFragBitInfo(16'b0000000000111111),.bFragBitInfo(16'b0000000100000011),.B1I0(NET_146),.B1I1(NET_495),.B1I2(fpgaio_out_dup_0[51]),.B1I3(fpgaio_oe_dup_0[51]),.T1I0(fpgaio_out_dup_0[51]),.T1I1(fpgaio_oe_dup_0[51]),.T1I2(NET_146),.T1I3(NET_495),.TB1S(NET_133),.C1Z(NET_486),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_B16_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_76),.B2I1(NET_75_CAND5_TLSBL_2_tpGCLKBUF),.B2I2(fpgaio_oe_dup_0[5]),.B2I3(fpgaio_out_dup_0[37]),.T2I0(NET_75_CAND5_TLSBL_2_tpGCLKBUF),.T2I1(fpgaio_out_dup_0[33]),.T2I2(fpgaio_oe_dup_0[1]),.T2I3(NET_76),.TB2S(GND),.B2Z(NET_827),.C2Z(NET_14),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_B16_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(fpgaio_oe_dup_0[27]),.T3I1(NET_72),.T3I2(fpgaio_oe_dup_0[59]),.T3I3(NET_75_CAND5_TLSBL_2_tpGCLKBUF),.C3Z(NET_684),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_B17_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_oe_dup_0[48]),.B0I1(NET_75),.B0I2(NET_72),.B0I3(fpgaio_oe_dup_0[16]),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.T0I0(NET_73),.T0I1(fpgaio_out_dup_0[16]),.T0I2(fpgaio_out_dup_0[48]),.T0I3(NET_76),.TB0S(GND),.B0Z(NET_429),.C0Z(NET_428),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_B17_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.T1I0(NET_72),.T1I1(NET_75),.T1I2(fpgaio_oe_dup_0[30]),.T1I3(fpgaio_oe_dup_0[62]),.C1Z(NET_756),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_B17_2 (.tFragBitInfo(16'b0101000011110000),.bFragBitInfo(16'b0001000000110000),.B2I0(fpgaio_oe_dup_0[41]),.B2I1(fpgaio_out_dup_0[9]),.B2I2(NET_239),.B2I3(NET_72),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_oe_dup_0[41]),.T2I1(fpgaio_out_dup_0[9]),.T2I2(NET_239),.T2I3(NET_72),.TB2S(NET_73),.C2Z(NET_240),.Q2Z(fpgaio_oe_dup_0[64]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_B17_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.T3I0(NET_73),.T3I1(NET_76),.T3I2(fpgaio_out_dup_0[25]),.T3I3(fpgaio_out_dup_0[57]),.C3Z(NET_641),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_B18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_147),.B0I1(fpgaio_oe_dup_0[44]),.B0I2(fpgaio_oe_dup_0[76]),.B0I3(NET_146),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B0Z(NET_308),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B18_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.T1I0(NET_147),.T1I1(fpgaio_oe_dup_0[38]),.T1I2(fpgaio_oe_dup_0[70]),.T1I3(NET_146),.C1Z(NET_794),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_B18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[76]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[70]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[62]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[38]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[48]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx4939z1_CAND3_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[47]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[47]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[41]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[51]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx4939z1_CAND3_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[32]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx4939z1_CAND3_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[35]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[33]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[59]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[46]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[60]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx4939z1_CAND3_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[62]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx4939z1_CAND3_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[37]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx4939z1_CAND3_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[33]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx4939z1_CAND3_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[51]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx4939z1_CAND3_BLSTL_2_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_2_padClk),.QRT(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[38]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_B25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_B25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_B25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_B25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx4939z1),.QCK(CLK_int_0__CAND0_BLSBL_2_padClk),.QRT(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[48]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[27]),.Q1EN(nx39840z1_CAND4_TLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx44608z1),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_3_padClk),.QRT(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx44608z1_CAND2_TLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C13_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_114),.B0I1(NET_143),.B0I2(fpgaio_in_int[21]),.B0I3(fpgaio_in_int[53]),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.T0I0(NET_114),.T0I1(NET_143),.T0I2(fpgaio_in_int[54]),.T0I3(fpgaio_in_int[22]),.TB0S(GND),.B0Z(NET_540),.C0Z(NET_563),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_C13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx39840z1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C13_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.T3I0(NET_114),.T3I1(NET_143),.T3I2(fpgaio_in_int[23]),.T3I3(fpgaio_in_int[55]),.TB3S(GND),.C3Z(NET_582),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_C14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_GNT_dup_0),.Q2EN(not_apb_fsm_1),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.Q2Z(lint_VALID_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx44608z1_CAND2_TLSBL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_3_padClk),.QRT(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_out_dup_0[59]),.B0I1(fpgaio_out_dup_0[27]),.B0I2(NET_76),.B0I3(NET_73_CAND3_TLSBL_3_tpGCLKBUF),.B0Z(NET_683),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C16_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(fpgaio_oe_dup_0[46]),.T1I1(fpgaio_oe_dup_0[14]),.T1I2(NET_72),.T1I3(NET_75_CAND5_TLSBL_3_tpGCLKBUF),.TB1S(GND),.C1Z(NET_356),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_C16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(fpgaio_oe_dup_0[32]),.B0I1(NET_147),.B0I2(NET_146),.B0I3(fpgaio_oe_dup_0[64]),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B0Z(NET_98),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[66]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(fpgaio_oe_dup_0[34]),.B2I1(NET_147),.B2I2(fpgaio_oe_dup_0[66]),.B2I3(NET_146),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B2Z(NET_896),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C17_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.T3I0(NET_76),.T3I1(fpgaio_out_dup_0[30]),.T3I2(NET_73),.T3I3(fpgaio_out_dup_0[62]),.C3Z(NET_755),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_C18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_146),.B0I1(NET_147),.B0I2(fpgaio_oe_dup_0[71]),.B0I3(fpgaio_oe_dup_0[39]),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B0Z(NET_594),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[71]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[68]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[72]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx9707z1_CAND5_BLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[39]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx9707z1_CAND5_BLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[34]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx9707z1_CAND5_BLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[43]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx9707z1_CAND5_BLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[32]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_C22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_C22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_C22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_C22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx4939z1_CAND3_BLSTL_3_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_3_padClk),.QRT(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[59]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D3_1 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx42928z2_CAND3_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p0_int[2]),.T1I1(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.T1I2(lint_WDATA_int[2]),.T1I3(GND),.TB1S(GND),.Q1Z(m0_oper0_wdata_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_D3_2 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42928z2_CAND3_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[3]),.T2I1(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.T2I2(GND),.T2I3(tcdm_rdata_p0_int[3]),.TB2S(GND),.Q2Z(m0_oper0_wdata_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_D3_3 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42928z2_CAND3_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p0_int[1]),.T3I1(lint_WDATA_int[1]),.T3I2(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper0_wdata_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_D4_0 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42928z2_CAND3_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[7]),.T0I1(tcdm_rdata_p0_int[7]),.T0I2(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.T0I3(GND),.TB0S(GND),.Q0Z(m0_oper0_wdata_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_D4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D4_3 (.tFragBitInfo(16'b0101010000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42928z2_CAND3_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.T3I2(tcdm_rdata_p0_int[9]),.T3I3(lint_WDATA_int[9]),.TB3S(GND),.Q3Z(m0_oper0_wdata_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_D7_0 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42928z2_CAND3_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[27]),.T0I1(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF),.T0I2(GND),.T0I3(tcdm_rdata_p0_int[27]),.TB0S(GND),.Q0Z(m0_oper0_wdata_dup_0[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_D7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_4_padClk),.QRT(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx44608z1_CAND2_TLSBL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D14_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_305),.B0I1(NET_307),.B0I2(NET_306),.B0I3(NET_304),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.T0I0(NET_305),.T0I1(NET_307),.T0I2(NET_306),.T0I3(NET_304),.TB0S(NET_308),.Q0Z(lint_RDATA_dup_0[12]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_D14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D15_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_94),.B0I1(NET_95),.B0I2(NET_96),.B0I3(NET_97),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.T0I0(NET_94),.T0I1(NET_95),.T0I2(NET_96),.T0I3(NET_97),.TB0S(NET_98),.Q0Z(lint_RDATA_dup_0[0]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_D15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D16_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.T0I0(NET_14),.T0I1(NET_12),.T0I2(NET_13),.T0I3(NET_11),.TB0S(GND),.Q0Z(lint_RDATA_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_D16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D16_2 (.tFragBitInfo(16'b0010000010100000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_73_CAND3_TLSBL_4_tpGCLKBUF),.B2I1(fpgaio_out_dup_0[14]),.B2I2(NET_55),.B2I3(fpgaio_oe_dup_0[78]),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.T2I0(NET_365),.T2I1(NET_76),.T2I2(NET_364),.T2I3(fpgaio_out_dup_0[46]),.TB2S(GND),.B2Z(NET_357),.C2Z(NET_355),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_D16_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_356),.B3I1(NET_354),.B3I2(NET_353),.B3I3(NET_355),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_4_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF),.T3I0(NET_353),.T3I1(NET_355),.T3I2(NET_356),.T3I3(NET_354),.TB3S(NET_357),.Q3Z(lint_RDATA_dup_0[14]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_D17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[78]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000100),.B2I0(GND),.B2I1(NET_55),.B2I2(GND),.B2I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B2Z(NET_147),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[65]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_oe_dup_0[75]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(fpgaio_oe_dup_0[75]),.B2I1(fpgaio_oe_dup_0[43]),.B2I2(NET_55),.B2I3(NET_72),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B2Z(NET_284),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[73]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx4939z1_CAND3_BLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[58]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_D20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_D20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx4939z1_CAND3_BLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[61]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_D20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx4939z1_CAND3_BLSTL_4_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[46]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_D20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_4_padClk),.QRT(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E1_0 (.tFragBitInfo(16'b1010110010100000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[7]),.T0I1(p0_cnt[5]),.T0I2(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T0I3(p0_fsm[3]),.TB0S(GND),.Q0Z(m0_oper0_waddr_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E1_1 (.tFragBitInfo(16'b1010101011000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[7]),.T1I1(p0_cnt[5]),.T1I2(p0_fsm[4]),.T1I3(NET_479),.TB1S(GND),.Q1Z(m0_oper0_raddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E1_2 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[0]),.T2I1(GND),.T2I2(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T2I3(GND),.TB2S(GND),.Q2Z(m0_oper0_waddr_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E1_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T3I1(lint_ADDR_int[1]),.T3I2(GND),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper0_waddr_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E2_0 (.tFragBitInfo(16'b1111100000001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T0I0(p0_fsm[4]),.T0I1(p0_cnt[9]),.T0I2(NET_479),.T0I3(lint_ADDR_int[11]),.TB0S(GND),.Q0Z(m0_oper0_raddr_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E2_1 (.tFragBitInfo(16'b1111100000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(p0_fsm[3]),.T1I1(p0_cnt[4]),.T1I2(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T1I3(lint_ADDR_int[6]),.TB1S(GND),.Q1Z(m0_oper0_waddr_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E2_2 (.tFragBitInfo(16'b1111100000001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T2I0(p0_fsm[3]),.T2I1(p0_cnt[9]),.T2I2(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T2I3(lint_ADDR_int[11]),.TB2S(GND),.Q2Z(m0_oper0_waddr_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E2_3 (.tFragBitInfo(16'b1111100000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(p0_fsm[4]),.T3I1(p0_cnt[4]),.T3I2(NET_479),.T3I3(lint_ADDR_int[6]),.TB3S(GND),.Q3Z(m0_oper0_raddr_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E3_0 (.tFragBitInfo(16'b1100101011000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T0I0(p0_fsm[3]),.T0I1(lint_ADDR_int[4]),.T0I2(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T0I3(p0_cnt[2]),.TB0S(GND),.Q0Z(m0_oper0_waddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E3_1 (.tFragBitInfo(16'b1111100000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(p0_cnt[1]),.T1I1(p0_fsm[3]),.T1I2(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T1I3(lint_ADDR_int[3]),.TB1S(GND),.Q1Z(m0_oper0_waddr_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E3_2 (.tFragBitInfo(16'b1110101001000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T2I0(NET_479),.T2I1(p0_fsm[4]),.T2I2(p0_cnt[1]),.T2I3(lint_ADDR_int[3]),.TB2S(GND),.Q2Z(m0_oper0_raddr_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E3_3 (.tFragBitInfo(16'b1110010010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(NET_479),.T3I1(p0_fsm[4]),.T3I2(lint_ADDR_int[4]),.T3I3(p0_cnt[2]),.TB3S(GND),.Q3Z(m0_oper0_raddr_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E4_2 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42928z2_CAND3_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[4]),.T2I1(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T2I2(GND),.T2I3(tcdm_rdata_p0_int[4]),.TB2S(GND),.Q2Z(m0_oper0_wdata_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E5_2 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42928z2_CAND3_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[19]),.T2I1(GND),.T2I2(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T2I3(tcdm_rdata_p0_int[19]),.TB2S(GND),.Q2Z(m0_oper0_wdata_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E5_3 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42928z2_CAND3_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p0_int[12]),.T3I1(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T3I2(lint_WDATA_int[12]),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper0_wdata_dup_0[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E6_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42928z2_CAND3_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[28]),.T3I1(tcdm_rdata_p0_int[28]),.T3I2(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper0_wdata_dup_0[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E7_0 (.tFragBitInfo(16'b0101000101000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42928z2_CAND3_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T0I2(lint_WDATA_int[25]),.T0I3(tcdm_rdata_p0_int[25]),.TB0S(GND),.Q0Z(m0_oper0_wdata_dup_0[25]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E7_3 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42928z2_CAND3_TLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_5_padClk),.QRT(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p0_int[23]),.T3I1(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF),.T3I2(lint_WDATA_int[23]),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper0_wdata_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx44608z1_CAND2_TLSBL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(m0_oper0_rmode_dup_0[0]),.B0I1(NET_143),.B0I2(fpgaio_in_int[0]),.B0I3(NET_142),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.B0Z(NET_137),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E10_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_in_int[2]),.T1I1(NET_143),.T1I2(m0_oper0_wmode_dup_0[0]),.T1I3(NET_142),.C1Z(NET_912),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_E10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper0_rmode_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wmode_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E12_0 (.tFragBitInfo(16'b0011001000010000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0EN(nx10146z2),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.T0I0(apb_fsm[1]),.T0I1(GND),.T0I2(nx10146z1),.T0I3(not_apb_fsm_0),.TB0S(GND),.Q0Z(apb_fsm[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.Q0DI(GND),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E12_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.T1I0(apb_fsm[0]),.T1I1(GND),.T1I2(GND),.T1I3(GND),.C1Z(not_apb_fsm_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_E12_2 (.tFragBitInfo(16'b0000000000110010),.bFragBitInfo(16'b1111110111111100),.B2I0(lint_GNT_dup_0),.B2I1(apb_fsm[0]),.B2I2(apb_fsm[1]),.B2I3(lint_REQ_int),.CD2S(GND),.Q2DI(GND),.Q2EN(nx10146z2),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.T2I0(lint_WEN_int),.T2I1(apb_fsm[0]),.T2I2(apb_fsm[1]),.T2I3(GND),.TB2S(GND),.B2Z(nx10146z2),.Q2Z(apb_fsm[1]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E12_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.QST(GND),.T3I0(lint_WEN_int),.T3I1(apb_fsm[0]),.T3I2(GND),.T3I3(GND),.TB3S(GND),.C3Z(nx10146z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_E13_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_537),.B0I1(NET_542),.B0I2(NET_922),.B0I3(NET_531),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T0I0(NET_537),.T0I1(NET_542),.T0I2(NET_922),.T0I3(NET_531),.TB0S(NET_547),.Q0Z(lint_RDATA_dup_0[21]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E13_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T1I0(lint_ADDR_int[6]),.T1I1(NET_91),.T1I2(NET_81),.T1I3(GND),.TB1S(GND),.C1Z(nx39840z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_E13_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_460),.B2I1(NET_919),.B2I2(NET_471),.B2I3(NET_466),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T2I0(NET_460),.T2I1(NET_919),.T2I2(NET_471),.T2I3(NET_466),.TB2S(NET_478),.Q2Z(lint_RDATA_dup_0[18]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E13_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_591),.B3I1(NET_592),.B3I2(NET_590),.B3I3(NET_593),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T3I0(NET_590),.T3I1(NET_593),.T3I2(NET_591),.T3I3(NET_592),.TB3S(NET_594),.Q3Z(lint_RDATA_dup_0[7]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E14_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_792),.B0I1(NET_790),.B0I2(NET_791),.B0I3(NET_793),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T0I0(NET_792),.T0I1(NET_790),.T0I2(NET_791),.T0I3(NET_793),.TB0S(NET_794),.Q0Z(lint_RDATA_dup_0[6]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E14_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B1I0(NET_584),.B1I1(NET_579),.B1I2(NET_923),.B1I3(NET_573),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T1I0(NET_923),.T1I1(NET_573),.T1I2(NET_584),.T1I3(NET_579),.TB1S(NET_589),.Q1Z(lint_RDATA_dup_0[23]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B2I0(apb_fsm[1]),.B2I1(GND),.B2I2(GND),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.B2Z(not_apb_fsm_1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E14_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_893),.B3I1(NET_894),.B3I2(NET_892),.B3I3(NET_895),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T3I0(NET_892),.T3I1(NET_895),.T3I2(NET_893),.T3I3(NET_894),.TB3S(NET_896),.Q3Z(lint_RDATA_dup_0[2]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_570),.B0I1(NET_81),.B0I2(NET_10),.B0I3(NET_673),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T0I0(NET_570),.T0I1(NET_81),.T0I2(NET_10),.T0I3(NET_673),.TB0S(lint_ADDR_int[4]),.C0Z(nx44608z1),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E15_1 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T1I0(lint_ADDR_int[5]),.T1I1(lint_ADDR_int[3]),.T1I2(lint_ADDR_int[6]),.T1I3(GND),.C1Z(NET_673),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_E15_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T2I0(NET_721),.T2I1(NET_719),.T2I2(NET_718),.T2I3(NET_720),.TB2S(GND),.Q2Z(lint_RDATA_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E15_3 (.tFragBitInfo(16'b0100110000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_5_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF),.T3I0(fpgaio_out_dup_0[61]),.T3I1(NET_730),.T3I2(NET_133),.T3I3(NET_729),.C3Z(NET_718),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_E16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_10),.B2I1(NET_570),.B2I2(lint_ADDR_int[2]),.B2I3(NET_673),.T2I0(NET_10),.T2I1(NET_570),.T2I2(lint_ADDR_int[2]),.T2I3(NET_673),.TB2S(lint_ADDR_int[4]),.C2Z(nx9707z1),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_E16_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_142),.T3I1(NET_143),.T3I2(fpgaio_in_int[12]),.T3I3(m0_oper0_wdsel_dup_0),.TB3S(GND),.C3Z(NET_324),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_E17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[67]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[79]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000000000000),.B0I0(lint_ADDR_int[5]),.B0I1(lint_ADDR_int[2]),.B0I2(NET_91),.B0I3(lint_ADDR_int[6]),.B0Z(nx4939z1),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000100000),.B2I0(lint_ADDR_int[5]),.B2I1(lint_ADDR_int[2]),.B2I2(NET_91),.B2I3(lint_ADDR_int[6]),.B2Z(nx19726z1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E20_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(NET_142),.T1I1(fpgaio_in_int[60]),.T1I2(m0_ram_control[28]),.T1I3(NET_114),.C1Z(NET_701),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_E20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(m0_ram_control[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper0_wdsel_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[20]),.Q2EN(nx9707z1_CAND5_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_oe_dup_0[52]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx4939z1_CAND3_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[60]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E22_0 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx12783z2_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T0I0(nx22245z2_CAND2_BLSTL_5_tpGCLKBUF),.T0I1(lint_WDATA_int[12]),.T0I2(GND),.T0I3(tcdm_rdata_p2_int[12]),.TB0S(GND),.Q0Z(m1_oper0_wdata_dup_0[12]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E22_3 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx12783z2_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T3I0(nx22245z2_CAND2_BLSTL_5_tpGCLKBUF),.T3I1(lint_WDATA_int[0]),.T3I2(tcdm_rdata_p2_int[0]),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper0_wdata_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E23_1 (.tFragBitInfo(16'b0101000101000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx12783z2_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(nx22245z2_CAND2_BLSTL_5_tpGCLKBUF),.T1I2(lint_WDATA_int[7]),.T1I3(tcdm_rdata_p2_int[7]),.TB1S(GND),.Q1Z(m1_oper0_wdata_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E23_2 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T2I0(nx22245z2_CAND2_BLSTL_5_tpGCLKBUF),.T2I1(tcdm_rdata_p2_int[10]),.T2I2(lint_WDATA_int[10]),.T2I3(GND),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_E24_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx12783z2_CAND4_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p2_int[15]),.T1I1(lint_WDATA_int[15]),.T1I2(nx22245z2_CAND2_BLSTL_5_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(m1_oper0_wdata_dup_0[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx4939z1_CAND3_BLSTL_5_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[56]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_5_padClk),.QRT(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E26_0 (.tFragBitInfo(16'b0000001100000010),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T0I0(nx22245z2_CAND2_BLSBL_5_tpGCLKBUF),.T0I1(GND),.T0I2(GND),.T0I3(p2_fsm[3]),.TB0S(GND),.C0Z(nx12783z2),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E26_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p2_int[18]),.T1I1(lint_WDATA_int[18]),.T1I2(nx22245z2_CAND2_BLSBL_5_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(m1_oper0_wdata_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E26_2 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[30]),.T2I1(tcdm_rdata_p2_int[30]),.T2I2(nx22245z2_CAND2_BLSBL_5_tpGCLKBUF),.T2I3(GND),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[30]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_E28_0 (.tFragBitInfo(16'b1110110000100000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T0I0(p2_cnt[3]),.T0I1(nx22245z2_CAND2_BLSBL_5_tpGCLKBUF),.T0I2(p2_fsm[3]),.T0I3(lint_ADDR_int[5]),.TB0S(GND),.Q0Z(m1_oper0_waddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_E28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_E28_3 (.tFragBitInfo(16'b1100110010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T3I0(p2_cnt[0]),.T3I1(lint_ADDR_int[2]),.T3I2(p2_fsm[3]),.T3I3(nx22245z2_CAND2_BLSBL_5_tpGCLKBUF),.TB3S(GND),.Q3Z(m1_oper0_waddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E29_0 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T0I0(nx22245z2_CAND2_BLSBL_5_tpGCLKBUF),.T0I1(GND),.T0I2(GND),.T0I3(lint_ADDR_int[1]),.TB0S(GND),.Q0Z(m1_oper0_waddr_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E29_1 (.tFragBitInfo(16'b1110110000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T1I0(p2_fsm[3]),.T1I1(nx22245z2_CAND2_BLSBL_5_tpGCLKBUF),.T1I2(p2_cnt[4]),.T1I3(lint_ADDR_int[6]),.TB1S(GND),.Q1Z(m1_oper0_waddr_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E29_2 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T2I0(nx22245z2_CAND2_BLSBL_5_tpGCLKBUF),.T2I1(lint_ADDR_int[0]),.T2I2(GND),.T2I3(GND),.TB2S(GND),.Q2Z(m1_oper0_waddr_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_E29_3 (.tFragBitInfo(16'b1110110000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T3I0(p2_fsm[3]),.T3I1(nx22245z2_CAND2_BLSBL_5_tpGCLKBUF),.T3I2(p2_cnt[1]),.T3I3(lint_ADDR_int[3]),.TB3S(GND),.Q3Z(m1_oper0_waddr_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E30_0 (.tFragBitInfo(16'b1110010010100000),.bFragBitInfo(16'b0001001100100000),.B0I0(NET_485),.B0I1(GND),.B0I2(m1_oper0_raddr_dup_0[6]),.B0I3(m1_oper0_raddr_dup_0[7]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx46309z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T0I0(NET_482_CAND3_BLSBL_5_tpGCLKBUF),.T0I1(NET_612),.T0I2(lint_ADDR_int[7]),.T0I3(p2_fsm_4__CAND5_BLSBL_5_tpGCLKBUF),.TB0S(GND),.B0Z(NET_612),.Q0Z(m1_oper0_raddr_dup_0[7]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E30_1 (.tFragBitInfo(16'b1000110110001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx46309z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T1I0(NET_482_CAND3_BLSBL_5_tpGCLKBUF),.T1I1(lint_ADDR_int[10]),.T1I2(NET_506),.T1I3(p2_fsm_4__CAND5_BLSBL_5_tpGCLKBUF),.TB1S(GND),.Q1Z(m1_oper0_raddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E30_2 (.tFragBitInfo(16'b0010000100000011),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T2I0(m1_oper0_raddr_dup_0[9]),.T2I1(GND),.T2I2(m1_oper0_raddr_dup_0[10]),.T2I3(NET_484),.TB2S(GND),.C2Z(NET_506),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_E30_3 (.tFragBitInfo(16'b1110001011000000),.bFragBitInfo(16'b1010101000001100),.B3I0(lint_ADDR_int[6]),.B3I1(p2_fsm_4__CAND5_BLSBL_5_tpGCLKBUF),.B3I2(NET_485),.B3I3(NET_482_CAND3_BLSBL_5_tpGCLKBUF),.CD3S(GND),.Q3DI(GND),.Q3EN(nx46309z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T3I0(NET_485),.T3I1(NET_482_CAND3_BLSBL_5_tpGCLKBUF),.T3I2(lint_ADDR_int[6]),.T3I3(p2_fsm_4__CAND5_BLSBL_5_tpGCLKBUF),.TB3S(m1_oper0_raddr_dup_0[6]),.Q3Z(m1_oper0_raddr_dup_0[6]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_E31_0 (.tFragBitInfo(16'b1010110010100000),.bFragBitInfo(16'b0111111110000000),.B0I0(m1_oper0_raddr_dup_0[7]),.B0I1(NET_485),.B0I2(m1_oper0_raddr_dup_0[6]),.B0I3(m1_oper0_raddr_dup_0[8]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx46309z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[8]),.T0I1(NET_569),.T0I2(NET_482_CAND3_BLSBL_5_tpGCLKBUF),.T0I3(p2_fsm_4__CAND5_BLSBL_5_tpGCLKBUF),.TB0S(GND),.B0Z(NET_569),.Q0Z(m1_oper0_raddr_dup_0[8]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_E31_1 (.tFragBitInfo(16'b1011100010001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx46309z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[11]),.T1I1(NET_482_CAND3_BLSBL_5_tpGCLKBUF),.T1I2(NET_483),.T1I3(p2_fsm_4__CAND5_BLSBL_5_tpGCLKBUF),.TB1S(GND),.Q1Z(m1_oper0_raddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_E31_2 (.tFragBitInfo(16'b0111100011110000),.bFragBitInfo(16'b1000000000000000),.B2I0(m1_oper0_raddr_dup_0[7]),.B2I1(NET_485),.B2I2(m1_oper0_raddr_dup_0[6]),.B2I3(m1_oper0_raddr_dup_0[8]),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T2I0(m1_oper0_raddr_dup_0[10]),.T2I1(NET_484),.T2I2(m1_oper0_raddr_dup_0[11]),.T2I3(m1_oper0_raddr_dup_0[9]),.TB2S(GND),.B2Z(NET_484),.C2Z(NET_483),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_E31_3 (.tFragBitInfo(16'b1010110010100000),.bFragBitInfo(16'b1010000011100100),.B3I0(NET_482_CAND3_BLSBL_5_tpGCLKBUF),.B3I1(p2_fsm_4__CAND5_BLSBL_5_tpGCLKBUF),.B3I2(lint_ADDR_int[9]),.B3I3(NET_484),.CD3S(GND),.Q3DI(GND),.Q3EN(nx46309z2),.QCK(CLK_int_0__CAND0_BLSBL_5_padClk),.QRT(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[9]),.T3I1(NET_484),.T3I2(NET_482_CAND3_BLSBL_5_tpGCLKBUF),.T3I3(p2_fsm_4__CAND5_BLSBL_5_tpGCLKBUF),.TB3S(m1_oper0_raddr_dup_0[9]),.Q3Z(m1_oper0_raddr_dup_0[9]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F1_0 (.tFragBitInfo(16'b1010110010100000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[10]),.T0I1(p0_cnt[8]),.T0I2(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T0I3(p0_fsm[3]),.TB0S(GND),.Q0Z(m0_oper0_waddr_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F1_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[0]),.T1I1(GND),.T1I2(NET_479),.T1I3(GND),.TB1S(GND),.Q1Z(m0_oper0_raddr_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_F1_2 (.tFragBitInfo(16'b1010101011000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[10]),.T2I1(p0_cnt[8]),.T2I2(p0_fsm[4]),.T2I3(NET_479),.TB2S(GND),.Q2Z(m0_oper0_raddr_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F1_3 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(lint_ADDR_int[1]),.T3I2(NET_479),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper0_raddr_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F2_0 (.tFragBitInfo(16'b1111000010001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T0I0(p0_fsm[4]),.T0I1(p0_cnt[7]),.T0I2(lint_ADDR_int[9]),.T0I3(NET_479),.TB0S(GND),.Q0Z(m0_oper0_raddr_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F2_1 (.tFragBitInfo(16'b1100110010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(p0_cnt[6]),.T1I1(lint_ADDR_int[8]),.T1I2(p0_fsm[4]),.T1I3(NET_479),.TB1S(GND),.Q1Z(m0_oper0_raddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_F2_2 (.tFragBitInfo(16'b1010101011000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[9]),.T2I1(p0_cnt[7]),.T2I2(p0_fsm[3]),.T2I3(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.TB2S(GND),.Q2Z(m0_oper0_waddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F2_3 (.tFragBitInfo(16'b1100110010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(p0_cnt[6]),.T3I1(lint_ADDR_int[8]),.T3I2(p0_fsm[3]),.T3I3(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.TB3S(GND),.Q3Z(m0_oper0_waddr_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F3_0 (.tFragBitInfo(16'b1101100010001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T0I0(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T0I1(lint_ADDR_int[5]),.T0I2(p0_cnt[3]),.T0I3(p0_fsm[3]),.TB0S(GND),.Q0Z(m0_oper0_waddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F3_1 (.tFragBitInfo(16'b1101100010001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx13379z2),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T1I1(lint_ADDR_int[2]),.T1I2(p0_cnt[0]),.T1I3(p0_fsm[3]),.TB1S(GND),.Q1Z(m0_oper0_waddr_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_F3_2 (.tFragBitInfo(16'b1101100010001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(NET_479),.T2I1(lint_ADDR_int[5]),.T2I2(p0_cnt[3]),.T2I3(p0_fsm[4]),.TB2S(GND),.Q2Z(m0_oper0_raddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F3_3 (.tFragBitInfo(16'b1100110010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx34850z5),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(p0_fsm[4]),.T3I1(lint_ADDR_int[2]),.T3I2(p0_cnt[0]),.T3I3(NET_479),.TB3S(GND),.Q3Z(m0_oper0_raddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F4_0 (.tFragBitInfo(16'b0000111000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42928z2_CAND3_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p0_int[26]),.T0I1(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T0I2(GND),.T0I3(lint_WDATA_int[26]),.TB0S(GND),.Q0Z(m0_oper0_wdata_dup_0[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F4_2 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42928z2_CAND3_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[10]),.T2I1(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T2I2(GND),.T2I3(tcdm_rdata_p0_int[10]),.TB2S(GND),.Q2Z(m0_oper0_wdata_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F5_1 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx42928z2_CAND3_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[15]),.T1I1(tcdm_rdata_p0_int[15]),.T1I2(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(m0_oper0_wdata_dup_0[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_F5_2 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42928z2_CAND3_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[11]),.T2I1(GND),.T2I2(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T2I3(tcdm_rdata_p0_int[11]),.TB2S(GND),.Q2Z(m0_oper0_wdata_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F5_3 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42928z2_CAND3_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p0_int[5]),.T3I1(lint_WDATA_int[5]),.T3I2(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper0_wdata_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F6_0 (.tFragBitInfo(16'b0101000101000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42928z2_CAND3_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T0I2(lint_WDATA_int[16]),.T0I3(tcdm_rdata_p0_int[16]),.TB0S(GND),.Q0Z(m0_oper0_wdata_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F6_3 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42928z2_CAND3_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p0_int[17]),.T3I1(lint_WDATA_int[17]),.T3I2(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper0_wdata_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F7_2 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42928z2_CAND3_TLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[31]),.T2I1(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF),.T2I2(GND),.T2I3(tcdm_rdata_p0_int[31]),.TB2S(GND),.Q2Z(m0_oper0_wdata_dup_0[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_6_padClk),.QRT(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F9_0 (.tFragBitInfo(16'b0100110001011111),.bFragBitInfo(16'b0100110000000000),.B0I0(fpgaio_oe_dup_0[11]),.B0I1(NET_929),.B0I2(NET_75_CAND5_TLSBL_6_tpGCLKBUF),.B0I3(apb_fsm[0]),.T0I0(fpgaio_oe_dup_0[11]),.T0I1(NET_929),.T0I2(NET_75_CAND5_TLSBL_6_tpGCLKBUF),.T0I3(apb_fsm[0]),.TB0S(lint_ADDR_int_11__CAND4_TLSBL_6_tpGCLKBUF),.C0Z(NET_930),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_F9_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(fpgaio_oe_dup_0[17]),.T1I1(lint_ADDR_int_11__CAND4_TLSBL_6_tpGCLKBUF),.T1I2(NET_75_CAND5_TLSBL_6_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.C1Z(NET_451),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_F9_2 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'b0000000000000000),.T2I0(fpgaio_oe_dup_0[19]),.T2I1(lint_ADDR_int_11__CAND4_TLSBL_6_tpGCLKBUF),.T2I2(NET_75_CAND5_TLSBL_6_tpGCLKBUF),.T2I3(GND),.TB2S(GND),.C2Z(NET_499),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_F9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B0I0(lint_REQ_int),.B0I1(GND),.B0I2(lint_GNT_dup_0),.B0I3(nx10146z1),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.QST(GND),.B0Z(nx7012z1),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F12_1 (.tFragBitInfo(16'b0000000000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.QST(GND),.T1I0(apb_fsm[0]),.T1I1(GND),.T1I2(GND),.T1I3(apb_fsm[1]),.C1Z(NET_10),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_F12_2 (.tFragBitInfo(16'b0000101000001100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2EN(nx7012z2),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.QST(GND),.T2I0(apb_fsm[0]),.T2I1(nx7012z1),.T2I2(GND),.T2I3(apb_fsm[1]),.TB2S(GND),.Q2Z(lint_GNT_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.Q2DI(GND),.T2CO());

	LOGIC_3 QL_INST_F12_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b0000000000000000),.B3I0(lint_GNT_dup_0),.B3I1(apb_fsm[0]),.B3I2(lint_REQ_int),.B3I3(lint_WEN_int),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(lint_REQ_int),.T3I1(lint_WEN_int),.T3I2(lint_GNT_dup_0),.T3I3(apb_fsm[0]),.TB3S(apb_fsm[1]),.C3Z(NET_79),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_F13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001101),.B0I0(apb_fsm[1]),.B0I1(apb_fsm[0]),.B0I2(GND),.B0I3(GND),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.B0Z(nx7012z2),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F13_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_552),.B3I1(NET_551),.B3I2(NET_553),.B3I3(NET_554),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.T3I0(NET_553),.T3I1(NET_554),.T3I2(NET_552),.T3I3(NET_551),.TB3S(NET_555),.Q3Z(lint_RDATA_dup_0[22]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F14_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0100110000000000),.B0I0(fpgaio_out_dup_0[56]),.B0I1(NET_626),.B0I2(NET_133),.B0I3(NET_625),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.T0I0(NET_616),.T0I1(NET_615),.T0I2(NET_614),.T0I3(NET_617),.TB0S(GND),.B0Z(NET_614),.Q0Z(lint_RDATA_dup_0[24]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F14_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.T1I0(NET_57),.T1I1(NET_31),.T1I2(NET_33),.T1I3(GND),.TB1S(GND),.C1Z(NET_75),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_F14_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000000010000),.B2I0(GND),.B2I1(GND),.B2I2(lint_ADDR_int[6]),.B2I3(lint_ADDR_int[5]),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.T2I0(NET_57),.T2I1(NET_74),.T2I2(NET_33),.T2I3(GND),.TB2S(GND),.B2Z(NET_57),.C2Z(NET_73),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_F14_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0000000000000000),.B3I0(NET_33),.B3I1(lint_ADDR_int[5]),.B3I2(NET_74),.B3I3(lint_ADDR_int_11__CAND4_TLSBL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.T3I0(NET_74),.T3I1(lint_ADDR_int_11__CAND4_TLSBL_6_tpGCLKBUF),.T3I2(NET_33),.T3I3(lint_ADDR_int[5]),.TB3S(lint_ADDR_int[6]),.C3Z(NET_142),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_F15_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000100010001000),.B0I0(NET_664),.B0I1(NET_665),.B0I2(fpgaio_out_dup_0[58]),.B0I3(NET_133),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.T0I0(NET_654),.T0I1(NET_653),.T0I2(NET_655),.T0I3(NET_656),.TB0S(GND),.B0Z(NET_653),.Q0Z(lint_RDATA_dup_0[26]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F15_1 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.T1I0(NET_695),.T1I1(NET_696),.T1I2(NET_697),.T1I3(NET_698),.TB1S(GND),.Q1Z(lint_RDATA_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_F15_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0100110000000000),.B2I0(fpgaio_out_dup_0[60]),.B2I1(NET_707),.B2I2(NET_133),.B2I3(NET_706),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.T2I0(NET_74),.T2I1(NET_29),.T2I2(NET_57),.T2I3(GND),.TB2S(GND),.B2Z(NET_695),.C2Z(NET_76),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_F15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_6_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F16_1 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int_11__CAND4_TLSBL_6_tpGCLKBUF),.T1I1(NET_57),.T1I2(NET_31),.T1I3(NET_29),.C1Z(NET_146),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_F16_2 (.tFragBitInfo(16'b0000000000000100),.bFragBitInfo(16'b0000000000000000),.T2I0(GND),.T2I1(lint_ADDR_int[4]),.T2I2(GND),.T2I3(lint_ADDR_int[3]),.TB2S(GND),.C2Z(NET_31),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_F16_3 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int_11__CAND4_TLSBL_6_tpGCLKBUF),.T3I1(NET_57),.T3I2(NET_74),.T3I3(NET_29),.C3Z(NET_133),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_F17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_oe_dup_0[77]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_oe_dup_0[69]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F19_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(NET_142),.T1I1(fpgaio_in_int[56]),.T1I2(m0_ram_control[24]),.T1I3(NET_114),.C1Z(NET_620),.Q1Z(m0_ram_control[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_F19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F22_2 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2_CAND4_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p2_int[23]),.T2I1(nx22245z2_CAND2_BLSTL_6_tpGCLKBUF),.T2I2(lint_WDATA_int[23]),.T2I3(GND),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F23_2 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2_CAND4_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_WDATA_int[5]),.T2I2(nx22245z2_CAND2_BLSTL_6_tpGCLKBUF),.T2I3(tcdm_rdata_p2_int[5]),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F24_1 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx12783z2_CAND4_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T1I0(nx22245z2_CAND2_BLSTL_6_tpGCLKBUF),.T1I1(GND),.T1I2(lint_WDATA_int[3]),.T1I3(tcdm_rdata_p2_int[3]),.TB1S(GND),.Q1Z(m1_oper0_wdata_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_F24_2 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2_CAND4_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_WDATA_int[11]),.T2I2(nx22245z2_CAND2_BLSTL_6_tpGCLKBUF),.T2I3(tcdm_rdata_p2_int[11]),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F24_3 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx12783z2_CAND4_BLSTL_6_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_6_padClk),.QRT(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(lint_WDATA_int[25]),.T3I2(nx22245z2_CAND2_BLSTL_6_tpGCLKBUF),.T3I3(tcdm_rdata_p2_int[25]),.TB3S(GND),.Q3Z(m1_oper0_wdata_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F25_0 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[6]),.T0I1(tcdm_rdata_p2_int[6]),.T0I2(nx22245z2_CAND2_BLSBL_6_tpGCLKBUF),.T0I3(GND),.TB0S(GND),.Q0Z(m1_oper0_wdata_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F25_1 (.tFragBitInfo(16'b0101000101000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(nx22245z2_CAND2_BLSBL_6_tpGCLKBUF),.T1I2(lint_WDATA_int[21]),.T1I3(tcdm_rdata_p2_int[21]),.TB1S(GND),.Q1Z(m1_oper0_wdata_dup_0[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_F25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F26_2 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T2I0(nx22245z2_CAND2_BLSBL_6_tpGCLKBUF),.T2I1(GND),.T2I2(lint_WDATA_int[24]),.T2I3(tcdm_rdata_p2_int[24]),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F26_3 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p2_int[17]),.T3I1(nx22245z2_CAND2_BLSBL_6_tpGCLKBUF),.T3I2(lint_WDATA_int[17]),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper0_wdata_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F27_0 (.tFragBitInfo(16'b0000000000010010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(GND),.QST(GND),.T0I0(p2_cnt[1]),.T0I1(GND),.T0I2(p2_cnt[0]),.T0I3(p2_fsm_0__CAND4_BLSBL_6_tpGCLKBUF),.TB0S(GND),.Q0Z(p2_cnt[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F27_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(GND),.QST(GND),.T1I0(GND),.T1I1(GND),.T1I2(p2_cnt[0]),.T1I3(p2_fsm_0__CAND4_BLSBL_6_tpGCLKBUF),.TB1S(GND),.Q1Z(p2_cnt[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_F27_2 (.tFragBitInfo(16'b0000000001101100),.bFragBitInfo(16'b0000000000010000),.B2I0(GND),.B2I1(p2_cnt[2]),.B2I2(control_in_int[18]),.B2I3(GND),.CD2S(GND),.Q2DI(GND),.Q2EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(GND),.QST(GND),.T2I0(p2_cnt[1]),.T2I1(p2_cnt[2]),.T2I2(p2_cnt[0]),.T2I3(p2_fsm_0__CAND4_BLSBL_6_tpGCLKBUF),.TB2S(GND),.B2Z(NET_172),.Q2Z(p2_cnt[2]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F27_3 (.tFragBitInfo(16'b1010001011111011),.bFragBitInfo(16'b0000000000000000),.B3I0(p2_cnt[0]),.B3I1(control_in_int[17]),.B3I2(p2_cnt[1]),.B3I3(control_in_int[16]),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(GND),.QST(GND),.T3I0(p2_cnt[1]),.T3I1(control_in_int[16]),.T3I2(p2_cnt[0]),.T3I3(control_in_int[17]),.TB3S(NET_172),.C3Z(NET_171),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_F28_0 (.tFragBitInfo(16'b1011001010110010),.bFragBitInfo(16'b1011001011110011),.B0I0(NET_171),.B0I1(control_in_int[19]),.B0I2(p2_cnt[3]),.B0I3(control_in_int[18]),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(GND),.QST(GND),.T0I0(NET_171),.T0I1(control_in_int[19]),.T0I2(p2_cnt[3]),.T0I3(control_in_int[18]),.TB0S(p2_cnt[2]),.C0Z(NET_170),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F28_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(GND),.QST(GND),.T1I0(p2_cnt[2]),.T1I1(p2_cnt[3]),.T1I2(p2_cnt[1]),.T1I3(p2_cnt[0]),.C1Z(NET_210),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_F28_2 (.tFragBitInfo(16'b0010001000100010),.bFragBitInfo(16'b0001001000100010),.B2I0(p2_cnt[3]),.B2I1(p2_fsm_0__CAND4_BLSBL_6_tpGCLKBUF),.B2I2(p2_cnt[1]),.B2I3(p2_cnt[0]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(GND),.QST(GND),.T2I0(p2_cnt[3]),.T2I1(p2_fsm_0__CAND4_BLSBL_6_tpGCLKBUF),.T2I2(p2_cnt[1]),.T2I3(p2_cnt[0]),.TB2S(p2_cnt[2]),.Q2Z(p2_cnt[3]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F28_3 (.tFragBitInfo(16'b0000000100010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(GND),.QST(GND),.T3I0(GND),.T3I1(p2_fsm_0__CAND4_BLSBL_6_tpGCLKBUF),.T3I2(NET_210),.T3I3(p2_cnt[4]),.TB3S(GND),.Q3Z(p2_cnt[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F29_0 (.tFragBitInfo(16'b1010110010100000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[4]),.T0I1(p2_cnt[2]),.T0I2(nx22245z2_CAND2_BLSBL_6_tpGCLKBUF),.T0I3(p2_fsm[3]),.TB0S(GND),.Q0Z(m1_oper0_waddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_F29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F30_1 (.tFragBitInfo(16'b1010111000000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx46309z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T1I0(NET_482_CAND3_BLSBL_6_tpGCLKBUF),.T1I1(p2_fsm_4__CAND5_BLSBL_6_tpGCLKBUF),.T1I2(m1_oper0_raddr_dup_0[2]),.T1I3(lint_ADDR_int[2]),.TB1S(GND),.Q1Z(m1_oper0_raddr_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_F30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_F31_0 (.tFragBitInfo(16'b1110010010100000),.bFragBitInfo(16'b0000000001101010),.B0I0(m1_oper0_raddr_dup_0[4]),.B0I1(m1_oper0_raddr_dup_0[2]),.B0I2(m1_oper0_raddr_dup_0[3]),.B0I3(GND),.CD0S(GND),.Q0DI(GND),.Q0EN(nx46309z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T0I0(NET_482_CAND3_BLSBL_6_tpGCLKBUF),.T0I1(NET_672),.T0I2(lint_ADDR_int[4]),.T0I3(p2_fsm_4__CAND5_BLSBL_6_tpGCLKBUF),.TB0S(GND),.B0Z(NET_672),.Q0Z(m1_oper0_raddr_dup_0[4]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_F31_1 (.tFragBitInfo(16'b0110101010101010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T1I0(m1_oper0_raddr_dup_0[5]),.T1I1(m1_oper0_raddr_dup_0[2]),.T1I2(m1_oper0_raddr_dup_0[3]),.T1I3(m1_oper0_raddr_dup_0[4]),.TB1S(GND),.C1Z(NET_650),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_F31_2 (.tFragBitInfo(16'b1101100010001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx46309z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T2I0(NET_482_CAND3_BLSBL_6_tpGCLKBUF),.T2I1(lint_ADDR_int[5]),.T2I2(NET_650),.T2I3(p2_fsm_4__CAND5_BLSBL_6_tpGCLKBUF),.TB2S(GND),.Q2Z(m1_oper0_raddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_F31_3 (.tFragBitInfo(16'b1110010010100000),.bFragBitInfo(16'b1010000010101100),.B3I0(lint_ADDR_int[3]),.B3I1(p2_fsm_4__CAND5_BLSBL_6_tpGCLKBUF),.B3I2(NET_482_CAND3_BLSBL_6_tpGCLKBUF),.B3I3(m1_oper0_raddr_dup_0[2]),.CD3S(GND),.Q3DI(GND),.Q3EN(nx46309z2),.QCK(CLK_int_0__CAND0_BLSBL_6_padClk),.QRT(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF),.QST(GND),.T3I0(NET_482_CAND3_BLSBL_6_tpGCLKBUF),.T3I1(m1_oper0_raddr_dup_0[2]),.T3I2(lint_ADDR_int[3]),.T3I3(p2_fsm_4__CAND5_BLSBL_6_tpGCLKBUF),.TB3S(m1_oper0_raddr_dup_0[3]),.Q3Z(m1_oper0_raddr_dup_0[3]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_F32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_F32_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m1_oper0_raddr_dup_0[5]),.T1I1(m1_oper0_raddr_dup_0[4]),.T1I2(m1_oper0_raddr_dup_0[2]),.T1I3(m1_oper0_raddr_dup_0[3]),.TB1S(GND),.C1Z(NET_485),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_F32_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_F32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000000000000),.B0I0(NET_786),.B0I1(GND),.B0I2(p0_cnt[6]),.B0I3(p0_cnt[7]),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.B0Z(NET_813),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G2_1 (.tFragBitInfo(16'b0000000000010010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.T1I0(NET_786),.T1I1(p0_fsm_0__CAND5_TLSTL_7_tpGCLKBUF),.T1I2(p0_cnt[6]),.T1I3(GND),.TB1S(GND),.Q1Z(p0_cnt[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_G2_2 (.tFragBitInfo(16'b0000011000001010),.bFragBitInfo(16'b0000100000000000),.B2I0(p0_cnt[5]),.B2I1(NET_745),.B2I2(GND),.B2I3(p0_cnt[4]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.T2I0(p0_cnt[5]),.T2I1(NET_745),.T2I2(p0_fsm_0__CAND5_TLSTL_7_tpGCLKBUF),.T2I3(p0_cnt[4]),.TB2S(GND),.B2Z(NET_786),.Q2Z(p0_cnt[5]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_G2_3 (.tFragBitInfo(16'b0001001100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.T3I0(NET_786),.T3I1(p0_fsm_0__CAND5_TLSTL_7_tpGCLKBUF),.T3I2(p0_cnt[6]),.T3I3(p0_cnt[7]),.TB3S(GND),.Q3Z(p0_cnt[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_G3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(p0_cnt[2]),.B0I1(p0_cnt[0]),.B0I2(p0_cnt[1]),.B0I3(p0_cnt[3]),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.B0Z(NET_745),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G3_1 (.tFragBitInfo(16'b1000110010101111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.T1I0(p0_cnt[7]),.T1I1(p0_cnt[6]),.T1I2(control_in_int[23]),.T1I3(control_in_int[22]),.C1Z(NET_189),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G3_3 (.tFragBitInfo(16'b0000000000010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.T3I0(GND),.T3I1(NET_745),.T3I2(p0_cnt[4]),.T3I3(p0_fsm_0__CAND5_TLSTL_7_tpGCLKBUF),.TB3S(GND),.Q3Z(p0_cnt[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_G4_0 (.tFragBitInfo(16'b0000000001101010),.bFragBitInfo(16'b1101110100001101),.B0I0(p0_cnt[5]),.B0I1(control_in_int[21]),.B0I2(p0_cnt[6]),.B0I3(control_in_int[22]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.T0I0(p0_cnt[2]),.T0I1(p0_cnt[0]),.T0I2(p0_cnt[1]),.T0I3(p0_fsm_0__CAND5_TLSTL_7_tpGCLKBUF),.TB0S(GND),.B0Z(NET_190),.Q0Z(p0_cnt[2]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G4_1 (.tFragBitInfo(16'b1101000011011101),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.T1I0(p0_cnt[3]),.T1I1(control_in_int[19]),.T1I2(control_in_int[20]),.T1I3(p0_cnt[4]),.C1Z(NET_192),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G4_2 (.tFragBitInfo(16'b0000000000000110),.bFragBitInfo(16'b1011000010111011),.B2I0(p0_cnt[5]),.B2I1(control_in_int[21]),.B2I2(p0_cnt[4]),.B2I3(control_in_int[20]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.T2I0(p0_cnt[1]),.T2I1(p0_cnt[0]),.T2I2(GND),.T2I3(p0_fsm_0__CAND5_TLSTL_7_tpGCLKBUF),.TB2S(GND),.B2Z(NET_191),.Q2Z(p0_cnt[1]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_G4_3 (.tFragBitInfo(16'b0011101100000000),.bFragBitInfo(16'b1100000011001100),.B3I0(NET_192),.B3I1(NET_189),.B3I2(NET_191),.B3I3(NET_190),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(GND),.QST(GND),.T3I0(NET_191),.T3I1(NET_190),.T3I2(NET_192),.T3I3(NET_189),.TB3S(NET_193),.C3Z(NET_187),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_G5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000100000),.B0I0(NET_198),.B0I1(GND),.B0I2(NET_79),.B0I3(lint_ADDR_int[14]),.CD0S(VCC),.Q0DI(control_in_int[0]),.Q0EN(VCC),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.B0Z(NET_479),.Q0Z(last_control[0]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G5_1 (.tFragBitInfo(16'b1100111011001100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(NET_198),.T1I1(NET_480),.T1I2(lint_ADDR_int[14]),.T1I3(NET_79),.TB1S(GND),.C1Z(nx34850z5),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_G5_2 (.tFragBitInfo(16'b1100010010100000),.bFragBitInfo(16'b1111001011110000),.B2I0(NET_198),.B2I1(lint_ADDR_int[14]),.B2I2(NET_206),.B2I3(NET_10),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(p0_fsm[3]),.T2I1(launch_p0),.T2I2(m0_oper0_we_dup_0),.T2I3(p0_fsm_0__CAND5_TLSTL_7_tpGCLKBUF),.TB2S(GND),.B2Z(nx13379z2),.C2Z(NET_206),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_G5_3 (.tFragBitInfo(16'b0001000001010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.T3I0(last_control[0]),.T3I1(launch_p0),.T3I2(control_in_int[0]),.T3I3(p0_fsm_0__CAND5_TLSTL_7_tpGCLKBUF),.C3Z(nx50997z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G6_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx42928z2_CAND3_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p0_int[21]),.T1I1(lint_WDATA_int[21]),.T1I2(nx34006z2_CAND2_TLSTL_7_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(m0_oper0_wdata_dup_0[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_G6_2 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42928z2_CAND3_TLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p0_int[29]),.T2I1(GND),.T2I2(nx34006z2_CAND2_TLSTL_7_tpGCLKBUF),.T2I3(lint_WDATA_int[29]),.TB2S(GND),.Q2Z(m0_oper0_wdata_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_G6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_7_padClk),.QRT(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.Q1Z(m0_oper0_rmode_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wdsel_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G11_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(m1_ram_control[29]),.T1I1(NET_124),.T1I2(NET_130),.T1I3(m0_m0_dataout_int[29]),.C1Z(NET_731),.Q1Z(m1_oper1_wdsel_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G11_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_734),.B2I1(NET_733),.B2I2(NET_731),.B2I3(NET_732),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T2I0(NET_668),.T2I1(NET_666),.T2I2(NET_667),.T2I3(NET_669),.TB2S(GND),.B2Z(NET_721),.C2Z(NET_656),.Q2Z(m1_ram_control[29]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_G11_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_dataout_int[26]),.T3I1(NET_124),.T3I2(NET_130),.T3I3(m1_ram_control[26]),.C3Z(NET_666),.Q3Z(m1_ram_control[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_131),.B0I1(NET_125),.B0I2(m1_m1_control[28]),.B0I3(m1_m0_dataout_int[28]),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.B0Z(NET_711),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G12_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(m0_m0_dataout_int[28]),.T1I1(NET_130),.T1I2(NET_124),.T1I3(m1_ram_control[28]),.C1Z(NET_708),.Q1Z(m1_m1_control[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_709),.B2I1(NET_710),.B2I2(NET_708),.B2I3(NET_711),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.B2Z(NET_698),.Q2Z(m1_m1_control[28]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G12_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_dataout_int[29]),.T3I1(NET_125),.T3I2(m1_m1_control[29]),.T3I3(NET_131),.C3Z(NET_734),.Q3Z(m1_ram_control[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G13_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx19381z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T0I0(NET_131),.T0I1(m1_m0_clr_dup_0),.T0I2(NET_128),.T0I3(m1_m1_clr_dup_0),.TB0S(GND),.C0Z(NET_443),.Q0Z(m1_m0_control[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G13_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[21]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(NET_128),.T1I1(NET_130),.T1I2(m1_ram_control[21]),.T1I3(m1_m0_control[21]),.TB1S(GND),.C1Z(NET_544),.Q1Z(m1_ram_control[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_G13_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0101011111110111),.B2I0(NET_34),.B2I1(m0_oper1_wdsel_dup_0),.B2I2(lint_ADDR_int[2]),.B2I3(m1_oper1_wdsel_dup_0),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx19381z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T2I0(NET_34),.T2I1(m0_oper1_wdsel_dup_0),.T2I2(lint_ADDR_int[2]),.T2I3(m1_oper1_wdsel_dup_0),.TB2S(NET_35),.C2Z(NET_337),.Q2Z(m1_m0_clr_dup_0),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_G13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx12574z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_outsel_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_907),.B0I1(NET_906),.B0I2(NET_905),.B0I3(NET_908),.CD0S(VCC),.Q0DI(lint_WDATA_int[2]),.Q0EN(nx41096z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.B0Z(NET_894),.Q0Z(m1_m1_control[2]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G14_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx12574z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_control[2]),.T1I1(m1_oper0_wmode_dup_0[0]),.T1I2(NET_131),.T1I3(NET_130),.C1Z(NET_908),.Q1Z(m0_m0_tc_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_m0_outsel_dup_0[0]),.B2I1(NET_128),.B2I2(m0_m0_outsel_dup_0[0]),.B2I3(NET_129),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.B2Z(NET_120),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G14_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx12574z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_outsel_dup_0[2]),.T3I1(NET_128),.T3I2(m0_m0_outsel_dup_0[2]),.T3I3(NET_129),.C3Z(NET_905),.Q3Z(m0_m0_outsel_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(m1_oper0_rmode_dup_0[0]),.B0I1(NET_130),.B0I2(NET_131),.B0I3(m1_m1_control[0]),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.B0Z(NET_123),.Q0Z(m1_m1_control[26]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G15_1 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx41096z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[12]),.T1I1(NET_9),.T1I2(lint_ADDR_int[13]),.T1I3(lint_ADDR_int[15]),.C1Z(NET_198),.Q1Z(m1_m1_control[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_m1_control[26]),.B2I1(NET_125),.B2I2(NET_131),.B2I3(m1_m0_dataout_int[26]),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.B2Z(NET_669),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G15_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(NET_122),.T3I1(NET_121),.T3I2(NET_123),.T3I3(NET_120),.C3Z(NET_96),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G16_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx36875z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[7]),.T0I1(apb_fsm[0]),.T0I2(lint_ADDR_int[2]),.T0I3(lint_ADDR_int[8]),.TB0S(GND),.C0Z(NET_33),.Q0Z(m1_m0_outsel_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx36875z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_outsel_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G16_2 (.tFragBitInfo(16'b1101111111111111),.bFragBitInfo(16'b0101111101111111),.B2I0(NET_35),.B2I1(lint_ADDR_int[2]),.B2I2(NET_117),.B2I3(fpgaio_in_int[19]),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx36875z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.T2I0(NET_35),.T2I1(lint_ADDR_int[2]),.T2I2(NET_117),.T2I3(fpgaio_in_int[19]),.TB2S(fpgaio_in_int[51]),.C2Z(NET_501),.Q2Z(m1_m0_outsel_dup_0[4]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_G16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx36875z1),.QCK(CLK_int_0__CAND0_TLSBL_7_padClk),.QRT(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF),.QST(GND),.Q3Z(m1_m0_outsel_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000100000),.B0I0(NET_33),.B0I1(GND),.B0I2(NET_117),.B0I3(GND),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B0Z(NET_143),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G17_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(NET_29),.T1I1(GND),.T1I2(NET_117),.T1I3(GND),.C1Z(NET_114),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_G17_2 (.tFragBitInfo(16'b1111111101111111),.bFragBitInfo(16'b0011111101111111),.B2I0(fpgaio_in_int[17]),.B2I1(NET_35),.B2I2(NET_117),.B2I3(lint_ADDR_int[2]),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[17]),.T2I1(NET_35),.T2I2(NET_117),.T2I3(lint_ADDR_int[2]),.TB2S(fpgaio_in_int[49]),.C2Z(NET_453),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_G17_3 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'b0000000000000000),.B3I0(lint_ADDR_int[5]),.B3I1(lint_ADDR_int[4]),.B3I2(lint_ADDR_int[6]),.B3I3(lint_ADDR_int[11]),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx58292z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[6]),.T3I1(lint_ADDR_int[11]),.T3I2(lint_ADDR_int[5]),.T3I3(lint_ADDR_int[4]),.TB3S(lint_ADDR_int[3]),.C3Z(NET_117),.Q3Z(fpgaio_oe_dup_0[74]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_G18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G18_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0101111101110111),.B2I0(NET_34),.B2I1(m0_oper0_rmode_dup_0[1]),.B2I2(m1_oper0_rmode_dup_0[1]),.B2I3(lint_ADDR_int[2]),.T2I0(NET_34),.T2I1(m0_oper0_rmode_dup_0[1]),.T2I2(m1_oper0_rmode_dup_0[1]),.T2I3(lint_ADDR_int[2]),.TB2S(NET_35),.C2Z(NET_26),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_G18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100000000000),.B0I0(NET_91),.B0I1(lint_ADDR_int[5]),.B0I2(lint_ADDR_int[6]),.B0I3(lint_ADDR_int[2]),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B0Z(nx49871z1),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_rmode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_rmode_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wmode_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G22_2 (.tFragBitInfo(16'b0000111000000010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p2_int[31]),.T2I1(nx22245z2_CAND2_BLSTL_7_tpGCLKBUF),.T2I2(GND),.T2I3(lint_WDATA_int[31]),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_G22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G23_0 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx12783z2_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p2_int[2]),.T0I1(nx22245z2_CAND2_BLSTL_7_tpGCLKBUF),.T0I2(lint_WDATA_int[2]),.T0I3(GND),.TB0S(GND),.Q0Z(m1_oper0_wdata_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G23_1 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx12783z2_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(lint_WDATA_int[28]),.T1I2(nx22245z2_CAND2_BLSTL_7_tpGCLKBUF),.T1I3(tcdm_rdata_p2_int[28]),.TB1S(GND),.Q1Z(m1_oper0_wdata_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_G23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_G23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G24_0 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx12783z2_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(lint_WDATA_int[14]),.T0I2(nx22245z2_CAND2_BLSTL_7_tpGCLKBUF),.T0I3(tcdm_rdata_p2_int[14]),.TB0S(GND),.Q0Z(m1_oper0_wdata_dup_0[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G24_2 (.tFragBitInfo(16'b0101000101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2_CAND4_BLSTL_7_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(nx22245z2_CAND2_BLSTL_7_tpGCLKBUF),.T2I2(lint_WDATA_int[19]),.T2I3(tcdm_rdata_p2_int[19]),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_G24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_7_padClk),.QRT(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G25_0 (.tFragBitInfo(16'b0101000101000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(nx22245z2_CAND2_BLSBL_7_tpGCLKBUF),.T0I2(lint_WDATA_int[8]),.T0I3(tcdm_rdata_p2_int[8]),.TB0S(GND),.Q0Z(m1_oper0_wdata_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G25_2 (.tFragBitInfo(16'b0000110000001010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p2_int[13]),.T2I1(lint_WDATA_int[13]),.T2I2(GND),.T2I3(nx22245z2_CAND2_BLSBL_7_tpGCLKBUF),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_G25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_G26_2 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_WDATA_int[22]),.T2I2(nx22245z2_CAND2_BLSBL_7_tpGCLKBUF),.T2I3(tcdm_rdata_p2_int[22]),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_G26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_G28_0 (.tFragBitInfo(16'b0000000000000110),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(GND),.QST(GND),.T0I0(p2_cnt[6]),.T0I1(NET_209),.T0I2(p2_fsm_0__CAND4_BLSBL_7_tpGCLKBUF),.T0I3(GND),.TB0S(GND),.Q0Z(p2_cnt[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_G28_1 (.tFragBitInfo(16'b0000011100001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(GND),.QST(GND),.T1I0(NET_210),.T1I1(p2_cnt[4]),.T1I2(p2_fsm_0__CAND4_BLSBL_7_tpGCLKBUF),.T1I3(p2_cnt[5]),.TB1S(GND),.Q1Z(p2_cnt[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_G28_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b1000001001000001),.B2I0(control_in_int[21]),.B2I1(p2_cnt[4]),.B2I2(control_in_int[20]),.B2I3(p2_cnt[5]),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(GND),.QST(GND),.T2I0(NET_210),.T2I1(p2_cnt[4]),.T2I2(GND),.T2I3(p2_cnt[5]),.TB2S(GND),.B2Z(NET_169),.C2Z(NET_209),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_G28_3 (.tFragBitInfo(16'b1101111101000101),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(GND),.QST(GND),.T3I0(control_in_int[21]),.T3I1(p2_cnt[4]),.T3I2(control_in_int[20]),.T3I3(p2_cnt[5]),.C3Z(NET_168),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_G29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_G29_1 (.tFragBitInfo(16'b1110001011000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.T1I0(p2_cnt[9]),.T1I1(nx22245z2_CAND2_BLSBL_7_tpGCLKBUF),.T1I2(lint_ADDR_int[11]),.T1I3(p2_fsm[3]),.TB1S(GND),.Q1Z(m1_oper0_waddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_G29_2 (.tFragBitInfo(16'b1011100010001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[8]),.T2I1(nx22245z2_CAND2_BLSBL_7_tpGCLKBUF),.T2I2(p2_cnt[6]),.T2I3(p2_fsm[3]),.TB2S(GND),.Q2Z(m1_oper0_waddr_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_G29_3 (.tFragBitInfo(16'b1110001011000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_7_padClk),.QRT(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF),.QST(GND),.T3I0(p2_cnt[5]),.T3I1(nx22245z2_CAND2_BLSBL_7_tpGCLKBUF),.T3I2(lint_ADDR_int[7]),.T3I3(p2_fsm[3]),.TB3S(GND),.Q3Z(m1_oper0_waddr_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_H2_0 (.tFragBitInfo(16'b0000000000000110),.bFragBitInfo(16'b0000000000000001),.B0I0(p0_cnt[9]),.B0I1(p0_cnt[10]),.B0I2(p0_cnt[11]),.B0I3(p0_cnt[8]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(GND),.QST(GND),.T0I0(NET_817),.T0I1(p0_cnt[10]),.T0I2(GND),.T0I3(p0_fsm_0__CAND5_TLSTL_8_tpGCLKBUF),.TB0S(GND),.B0Z(NET_197),.Q0Z(p0_cnt[10]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H2_1 (.tFragBitInfo(16'b0000000001111000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(GND),.QST(GND),.T1I0(NET_817),.T1I1(p0_cnt[10]),.T1I2(p0_cnt[11]),.T1I3(p0_fsm_0__CAND5_TLSTL_8_tpGCLKBUF),.TB1S(GND),.Q1Z(p0_cnt[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H2_2 (.tFragBitInfo(16'b0000011000001010),.bFragBitInfo(16'b0000100000000000),.B2I0(p0_cnt[9]),.B2I1(NET_813),.B2I2(GND),.B2I3(p0_cnt[8]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(GND),.QST(GND),.T2I0(p0_cnt[9]),.T2I1(NET_813),.T2I2(p0_fsm_0__CAND5_TLSTL_8_tpGCLKBUF),.T2I3(p0_cnt[8]),.TB2S(GND),.B2Z(NET_817),.Q2Z(p0_cnt[9]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_H2_3 (.tFragBitInfo(16'b0000000100000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(GND),.QST(GND),.T3I0(GND),.T3I1(NET_813),.T3I2(p0_fsm_0__CAND5_TLSTL_8_tpGCLKBUF),.T3I3(p0_cnt[8]),.TB3S(GND),.Q3Z(p0_cnt[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_H3_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(GND),.QST(GND),.T0I0(p0_fsm_0__CAND5_TLSTL_8_tpGCLKBUF),.T0I1(GND),.T0I2(GND),.T0I3(p0_cnt[0]),.TB0S(GND),.Q0Z(p0_cnt[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H3_1 (.tFragBitInfo(16'b0101000001010000),.bFragBitInfo(16'b0000011000001010),.B1I0(p0_cnt[3]),.B1I1(p0_cnt[1]),.B1I2(p0_fsm_0__CAND5_TLSTL_8_tpGCLKBUF),.B1I3(p0_cnt[0]),.CD1S(GND),.Q1DI(GND),.Q1EN(nx48658z2),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(GND),.QST(GND),.T1I0(p0_fsm_0__CAND5_TLSTL_8_tpGCLKBUF),.T1I1(p0_cnt[0]),.T1I2(p0_cnt[3]),.T1I3(p0_cnt[1]),.TB1S(p0_cnt[2]),.Q1Z(p0_cnt[3]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(GND),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H3_3 (.tFragBitInfo(16'b0000101000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(GND),.QST(GND),.T3I0(NET_197),.T3I1(p0_cnt[7]),.T3I2(GND),.T3I3(control_in_int[23]),.C3Z(NET_188),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H4_0 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000011110010),.B0I0(control_in_int[16]),.B0I1(p0_cnt[0]),.B0I2(control_in_int[17]),.B0I3(p0_cnt[1]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42928z2_CAND3_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[6]),.T0I1(nx34006z2_CAND2_TLSTL_8_tpGCLKBUF),.T0I2(GND),.T0I3(tcdm_rdata_p0_int[6]),.TB0S(GND),.B0Z(NET_196),.Q0Z(m0_oper0_wdata_dup_0[6]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H4_1 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(p0_cnt[3]),.T1I2(GND),.T1I3(control_in_int[19]),.C1Z(NET_194),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_H4_2 (.tFragBitInfo(16'b0000101000001011),.bFragBitInfo(16'b0000000000000010),.B2I0(p0_cnt[2]),.B2I1(NET_196),.B2I2(NET_194),.B2I3(NET_195),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T2I0(p0_cnt[2]),.T2I1(NET_196),.T2I2(NET_194),.T2I3(NET_195),.TB2S(control_in_int[18]),.C2Z(NET_193),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_H4_3 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(control_in_int[16]),.T3I1(p0_cnt[0]),.T3I2(control_in_int[17]),.T3I3(GND),.C3Z(NET_195),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H5_0 (.tFragBitInfo(16'b0000001100000010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0EN(VCC),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(nx50997z2),.T0I1(GND),.T0I2(GND),.T0I3(nx50997z1),.TB0S(GND),.Q0Z(launch_p0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.Q0DI(GND),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H5_1 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx42928z2_CAND3_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T1I0(nx34006z2_CAND2_TLSTL_8_tpGCLKBUF),.T1I1(tcdm_rdata_p0_int[8]),.T1I2(lint_WDATA_int[8]),.T1I3(GND),.TB1S(GND),.Q1Z(m0_oper0_wdata_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H5_2 (.tFragBitInfo(16'b0000000000001110),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2EN(VCC),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T2I0(nx34006z2_CAND2_TLSTL_8_tpGCLKBUF),.T2I1(nx34006z1),.T2I2(GND),.T2I3(GND),.TB2S(GND),.Q2Z(m0_oper0_we_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.Q2DI(GND),.T2CO());

	LOGIC_3 QL_INST_H5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H6_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx42928z2_CAND3_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p0_int[18]),.T1I1(lint_WDATA_int[18]),.T1I2(nx34006z2_CAND2_TLSTL_8_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(m0_oper0_wdata_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H6_2 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42928z2_CAND3_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T2I0(nx34006z2_CAND2_TLSTL_8_tpGCLKBUF),.T2I1(lint_WDATA_int[14]),.T2I2(GND),.T2I3(tcdm_rdata_p0_int[14]),.TB2S(GND),.Q2Z(m0_oper0_wdata_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_H6_3 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(NET_198),.T3I1(lint_ADDR_int[14]),.T3I2(NET_10),.T3I3(GND),.C3Z(nx34006z2),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H7_0 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42928z2_CAND3_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(nx34006z2_CAND2_TLSTL_8_tpGCLKBUF),.T0I1(lint_WDATA_int[30]),.T0I2(tcdm_rdata_p0_int[30]),.T0I3(GND),.TB0S(GND),.Q0Z(m0_oper0_wdata_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H7_1 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx42928z2_CAND3_TLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.T1I0(nx34006z2_CAND2_TLSTL_8_tpGCLKBUF),.T1I1(GND),.T1I2(lint_WDATA_int[22]),.T1I3(tcdm_rdata_p0_int[22]),.TB1S(GND),.Q1Z(m0_oper0_wdata_dup_0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTL_8_padClk),.QRT(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H11_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T0I0(NET_129),.T0I1(NET_124),.T0I2(m0_m0_control[21]),.T0I3(m0_m0_dataout_int[21]),.TB0S(GND),.C0Z(NET_543),.Q0Z(m0_oper0_wmode_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H11_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[23]),.Q1EN(nx1800z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_129),.T1I1(NET_124),.T1I2(m0_m0_dataout_int[22]),.T1I3(m0_m0_control[22]),.TB1S(GND),.C1Z(NET_565),.Q1Z(m0_m0_control[23]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_H11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_129),.B2I1(m0_m0_dataout_int[23]),.B2I2(NET_124),.B2I3(m0_m0_control[23]),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx1800z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.B2Z(NET_585),.Q2Z(m0_m0_control[21]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx1800z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_control[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H12_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx19381z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T0I0(NET_128),.T0I1(m1_m0_sat_dup_0),.T0I2(m1_m1_sat_dup_0),.T0I3(NET_131),.TB0S(GND),.C0Z(NET_463),.Q0Z(m1_m0_sat_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H12_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx19381z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_125),.T1I1(m0_m0_dataout_int[18]),.T1I2(NET_124),.T1I3(m1_m0_dataout_int[18]),.TB1S(GND),.C1Z(NET_477),.Q1Z(m1_m0_control[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_H12_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T2I0(NET_565),.T2I1(NET_567),.T2I2(NET_566),.T2I3(NET_568),.TB2S(GND),.C2Z(NET_551),.Q2Z(m1_ram_control[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_H12_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T3I0(NET_128),.T3I1(NET_130),.T3I2(m1_ram_control[22]),.T3I3(m1_m0_control[22]),.C3Z(NET_566),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(m1_m0_control[23]),.B0I1(NET_130),.B0I2(m1_ram_control[23]),.B0I3(NET_128),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx19381z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.B0Z(NET_586),.Q0Z(m1_m0_control[23]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H13_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[21]),.Q1EN(nx32122z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_545),.T1I1(NET_544),.T1I2(NET_546),.T1I3(NET_543),.TB1S(GND),.C1Z(NET_547),.Q1Z(m1_m1_control[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_H13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[23]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.Q2Z(m1_ram_control[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H13_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx32122z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T3I0(NET_125),.T3I1(m1_m0_dataout_int[21]),.T3I2(m1_m1_control[21]),.T3I3(NET_131),.TB3S(GND),.C3Z(NET_546),.Q3Z(m1_m1_sat_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_H14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100000000000),.B0I0(NET_912),.B0I1(NET_911),.B0I2(GND),.B0I3(NET_910),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.B0Z(NET_895),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H14_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx36875z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_128),.T1I1(m0_m0_tc_dup_0),.T1I2(NET_129),.T1I3(m1_m0_tc_dup_0),.C1Z(NET_803),.Q1Z(m1_m0_control[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_H14_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_128),.B2I1(m0_m0_control[7]),.B2I2(m1_m0_control[7]),.B2I3(NET_129),.CD2S(VCC),.Q2DI(lint_WDATA_int[7]),.Q2EN(nx12574z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T2I0(NET_585),.T2I1(NET_586),.T2I2(NET_588),.T2I3(NET_587),.TB2S(GND),.B2Z(NET_603),.C2Z(NET_589),.Q2Z(m0_m0_control[7]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_H14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx12574z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_outsel_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(m1_m0_dataout_int[22]),.B0I1(NET_131),.B0I2(m1_m1_control[22]),.B0I3(NET_125),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx32122z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.B0Z(NET_568),.Q0Z(m1_m1_control[23]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H15_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[22]),.Q1EN(nx32122z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_125),.T1I1(NET_124),.T1I2(m1_m0_dataout_int[19]),.T1I3(m0_m0_dataout_int[19]),.TB1S(GND),.C1Z(NET_492),.Q1Z(m1_m1_control[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_H15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_125),.B2I1(NET_131),.B2I2(m1_m1_control[24]),.B2I3(m1_m0_dataout_int[24]),.CD2S(VCC),.Q2DI(lint_WDATA_int[24]),.Q2EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.B2Z(NET_630),.Q2Z(m1_m1_control[24]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H15_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx36875z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_dataout_int[23]),.T3I1(NET_131),.T3I2(NET_125),.T3I3(m1_m1_control[23]),.TB3S(GND),.C3Z(NET_588),.Q3Z(m1_m0_outsel_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_H16_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_28),.B0I1(NET_41),.B0I2(fpgaio_in_int[57]),.B0I3(m0_m0_dataout_int[25]),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(lint_ADDR_int[4]),.T0I2(lint_ADDR_int[3]),.T0I3(GND),.TB0S(GND),.B0Z(NET_639),.C0Z(NET_74),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H16_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_28),.T1I1(NET_41),.T1I2(m0_m0_dataout_int[27]),.T1I3(fpgaio_in_int[59]),.C1Z(NET_681),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_H16_2 (.tFragBitInfo(16'b0100110001001100),.bFragBitInfo(16'b0000000001001100),.B2I0(NET_27),.B2I1(NET_337),.B2I2(m0_m0_mode_dup_0[1]),.B2I3(fpgaio_in_int[45]),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx32122z1),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T2I0(NET_27),.T2I1(NET_337),.T2I2(m0_m0_mode_dup_0[1]),.T2I3(fpgaio_in_int[45]),.TB2S(NET_28),.C2Z(NET_333),.Q2Z(m1_m1_clr_dup_0),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_H16_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBL_8_padClk),.QRT(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF),.QST(GND),.T3I0(NET_28),.T3I1(NET_41),.T3I2(fpgaio_in_int[62]),.T3I3(m0_m0_dataout_int[30]),.C3Z(NET_753),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx36875z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_tc_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx36875z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_outsel_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[64]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H18_1 (.tFragBitInfo(16'b0000000000000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[7]),.T1I1(lint_ADDR_int[2]),.T1I2(apb_fsm[0]),.T1I3(lint_ADDR_int[8]),.TB1S(GND),.C1Z(NET_29),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_H18_2 (.tFragBitInfo(16'b0100010011001100),.bFragBitInfo(16'b0000010000001100),.B2I0(NET_27),.B2I1(NET_26),.B2I2(fpgaio_in_int[33]),.B2I3(m0_m0_outsel_dup_0[1]),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T2I0(NET_27),.T2I1(NET_26),.T2I2(fpgaio_in_int[33]),.T2I3(m0_m0_outsel_dup_0[1]),.TB2S(NET_28),.C2Z(NET_17),.Q2Z(fpgaio_out_dup_0[65]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_H18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[74]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[77]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H20_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(NET_114),.T3I1(NET_142),.T3I2(fpgaio_in_int[61]),.T3I3(m0_ram_control[29]),.C3Z(NET_724),.Q3Z(m0_ram_control[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_H21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[15]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.Q0Z(m0_ram_control[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H21_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T1I0(NET_27),.T1I1(NET_28),.T1I2(fpgaio_in_int[46]),.T1I3(m0_m0_osel_dup_0),.TB1S(GND),.C1Z(NET_371),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_H21_2 (.tFragBitInfo(16'b0111011100000000),.bFragBitInfo(16'b0000011100000000),.B2I0(NET_27),.B2I1(m0_m0_csel_dup_0),.B2I2(fpgaio_in_int[47]),.B2I3(NET_404),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T2I0(NET_27),.T2I1(m0_m0_csel_dup_0),.T2I2(fpgaio_in_int[47]),.T2I3(NET_404),.TB2S(NET_28),.C2Z(NET_401),.Q2Z(m1_ram_control[15]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_H21_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001101111111111),.B3I0(lint_ADDR_int[2]),.B3I1(m0_ram_control[15]),.B3I2(m1_ram_control[15]),.B3I3(NET_34),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(m1_ram_control[15]),.T3I1(NET_34),.T3I2(lint_ADDR_int[2]),.T3I3(m0_ram_control[15]),.TB3S(NET_35),.C3Z(NET_404),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_H22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H22_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx12783z2_CAND4_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[27]),.T3I1(tcdm_rdata_p2_int[27]),.T3I2(nx22245z2_CAND2_BLSTL_8_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper0_wdata_dup_0[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_H23_0 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx12783z2_CAND4_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[20]),.T0I1(tcdm_rdata_p2_int[20]),.T0I2(nx22245z2_CAND2_BLSTL_8_tpGCLKBUF),.T0I3(GND),.TB0S(GND),.Q0Z(m1_oper0_wdata_dup_0[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H24_1 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx12783z2_CAND4_BLSTL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p2_int[9]),.T1I1(nx22245z2_CAND2_BLSTL_8_tpGCLKBUF),.T1I2(lint_WDATA_int[9]),.T1I3(GND),.TB1S(GND),.Q1Z(m1_oper0_wdata_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_H24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_H24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTL_8_padClk),.QRT(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_H26_0 (.tFragBitInfo(16'b1111111100001000),.bFragBitInfo(16'b1111111111011000),.B0I0(p2_fsm_0__CAND4_BLSBL_8_tpGCLKBUF),.B0I1(launch_p2),.B0I2(p2_fsm_4__CAND5_BLSBL_8_tpGCLKBUF),.B0I3(NET_482_CAND3_BLSBL_8_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.T0I0(p2_fsm_0__CAND4_BLSBL_8_tpGCLKBUF),.T0I1(launch_p2),.T0I2(p2_fsm_4__CAND5_BLSBL_8_tpGCLKBUF),.T0I3(NET_482_CAND3_BLSBL_8_tpGCLKBUF),.TB0S(tcdm_req_p2_dup_0),.C0Z(nx46309z2),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H26_1 (.tFragBitInfo(16'b0000000001010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1EN(VCC),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(nx22245z2_CAND2_BLSBL_8_tpGCLKBUF),.T1I2(nx22245z1),.T1I3(GND),.TB1S(GND),.Q1Z(m1_oper0_we_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.Q1DI(GND),.T1CO());

	LOGIC_2 QL_INST_H26_2 (.tFragBitInfo(16'b0000000000001110),.bFragBitInfo(16'b0000001000001010),.B2I0(control_in_int[2]),.B2I1(launch_p2),.B2I2(last_control[2]),.B2I3(p2_fsm_0__CAND4_BLSBL_8_tpGCLKBUF),.CD2S(GND),.Q2EN(VCC),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.T2I0(nx50995z3),.T2I1(nx50995z1),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(nx50995z1),.Q2Z(launch_p2),.B2CO(),.C2Z(),.Q2DI(GND),.T2CO());

	LOGIC_3 QL_INST_H26_3 (.tFragBitInfo(16'b1111111100001000),.bFragBitInfo(16'b1111111011001110),.B3I0(p2_fsm[3]),.B3I1(nx22245z2_CAND2_BLSBL_8_tpGCLKBUF),.B3I2(p2_fsm_0__CAND4_BLSBL_8_tpGCLKBUF),.B3I3(launch_p2),.CD3S(VCC),.Q3DI(control_in_int[2]),.Q3EN(VCC),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.T3I0(p2_fsm_0__CAND4_BLSBL_8_tpGCLKBUF),.T3I1(launch_p2),.T3I2(p2_fsm[3]),.T3I3(nx22245z2_CAND2_BLSBL_8_tpGCLKBUF),.TB3S(m1_oper0_we_dup_0),.C3Z(nx22012z2),.Q3Z(last_control[2]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_H28_0 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b1011001010111011),.B0I0(p2_cnt[7]),.B0I1(control_in_int[23]),.B0I2(p2_cnt[6]),.B0I3(control_in_int[22]),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(GND),.QST(GND),.T0I0(GND),.T0I1(p2_cnt[7]),.T0I2(p2_cnt[6]),.T0I3(NET_209),.TB0S(GND),.B0Z(NET_166),.C0Z(NET_208),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_H28_1 (.tFragBitInfo(16'b0100110001000100),.bFragBitInfo(16'b1100111100000000),.B1I0(NET_169),.B1I1(NET_168),.B1I2(NET_167),.B1I3(NET_166),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(GND),.QST(GND),.T1I0(NET_167),.T1I1(NET_166),.T1I2(NET_169),.T1I3(NET_168),.TB1S(NET_170),.C1Z(NET_164),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_H28_2 (.tFragBitInfo(16'b0001001000100010),.bFragBitInfo(16'b1001000000001001),.B2I0(p2_cnt[7]),.B2I1(control_in_int[23]),.B2I2(p2_cnt[6]),.B2I3(control_in_int[22]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(GND),.QST(GND),.T2I0(p2_cnt[7]),.T2I1(p2_fsm_0__CAND4_BLSBL_8_tpGCLKBUF),.T2I2(p2_cnt[6]),.T2I3(NET_209),.TB2S(GND),.B2Z(NET_167),.Q2Z(p2_cnt[7]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_H28_3 (.tFragBitInfo(16'b0000000000010010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(GND),.QST(GND),.T3I0(NET_208),.T3I1(p2_fsm_0__CAND4_BLSBL_8_tpGCLKBUF),.T3I2(p2_cnt[8]),.T3I3(GND),.TB3S(GND),.Q3Z(p2_cnt[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_H29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_H29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_H29_2 (.tFragBitInfo(16'b1111100000001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.T2I0(p2_fsm[3]),.T2I1(p2_cnt[7]),.T2I2(nx22245z2_CAND2_BLSBL_8_tpGCLKBUF),.T2I3(lint_ADDR_int[9]),.TB2S(GND),.Q2Z(m1_oper0_waddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_H29_3 (.tFragBitInfo(16'b1100101011000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx22012z2),.QCK(CLK_int_0__CAND0_BLSBL_8_padClk),.QRT(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF),.QST(GND),.T3I0(p2_fsm[3]),.T3I1(lint_ADDR_int[10]),.T3I2(nx22245z2_CAND2_BLSBL_8_tpGCLKBUF),.T3I3(p2_cnt[8]),.TB3S(GND),.Q3Z(m1_oper0_waddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_I3_0 (.tFragBitInfo(16'b0000010000000100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0EN(nx18527z1),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.T0I0(not_tcdm_wen_p0),.T0I1(nx21518z1),.T0I2(GND),.T0I3(GND),.TB0S(GND),.Q0Z(p0_fsm[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.Q0DI(GND),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I3_1 (.tFragBitInfo(16'b0011001000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx42928z2),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(nx34006z2),.T1I1(GND),.T1I2(tcdm_rdata_p0_int[0]),.T1I3(lint_WDATA_int[0]),.TB1S(GND),.Q1Z(m0_oper0_wdata_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_I3_2 (.tFragBitInfo(16'b1011101010101010),.bFragBitInfo(16'b0000000000000001),.B2I0(GND),.B2I1(tcdm_wen_p0_dup_0),.B2I2(GND),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.T2I0(p0_fsm[0]),.T2I1(NET_187),.T2I2(p0_fsm[4]),.T2I3(NET_188),.TB2S(GND),.B2Z(not_tcdm_wen_p0),.C2Z(nx21518z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001000),.B0I0(RESET_int[0]),.B0I1(NET_186),.B0I2(p0_fsm[4]),.B0I3(NET_217),.B0Z(nx48658z2),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I4_1 (.tFragBitInfo(16'b0000010011001100),.bFragBitInfo(16'b0111011100000000),.B1I0(p0_fsm[3]),.B1I1(NET_217),.B1I2(NET_188),.B1I3(NET_216),.T1I0(NET_188),.T1I1(NET_216),.T1I2(p0_fsm[3]),.T1I3(NET_217),.TB1S(NET_187),.C1Z(nx18527z1),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_I4_2 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(tcdm_wen_p0_dup_0),.T2I1(NET_187),.T2I2(p0_fsm[4]),.T2I3(NET_188),.TB2S(GND),.C2Z(nx20521z1),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_I4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I5_0 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b1111111100100000),.B0I0(NET_198),.B0I1(lint_ADDR_int[14]),.B0I2(NET_10),.B0I3(p0_fsm[3]),.T0I0(tcdm_wen_p0_dup_0),.T0I1(GND),.T0I2(p0_fsm[4]),.T0I3(tcdm_valid_p0_int_CAND3_TLSTR_9_tpGCLKBUF),.TB0S(GND),.B0Z(nx42928z2),.C0Z(nx34006z1),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_I5_1 (.tFragBitInfo(16'b1011101100001011),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(launch_p0),.T1I1(p0_fsm[0]),.T1I2(p0_fsm[4]),.T1I3(tcdm_valid_p0_int_CAND3_TLSTR_9_tpGCLKBUF),.TB1S(GND),.C1Z(NET_216),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_I5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I5_3 (.tFragBitInfo(16'b1010110000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(tcdm_req_p0_dup_0),.T3I1(p0_fsm[0]),.T3I2(p0_fsm[4]),.T3I3(launch_p0),.TB3S(GND),.C3Z(NET_480),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_I6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I6_2 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42928z2),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.T2I0(nx34006z2),.T2I1(GND),.T2I2(lint_WDATA_int[13]),.T2I3(tcdm_rdata_p0_int[13]),.TB2S(GND),.Q2Z(m0_oper0_wdata_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_I6_3 (.tFragBitInfo(16'b0011000000100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42928z2),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p0_int[20]),.T3I1(GND),.T3I2(lint_WDATA_int[20]),.T3I3(nx34006z2),.TB3S(GND),.Q3Z(m0_oper0_wdata_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_I7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[24]),.Q0EN(tcdm_valid_p0_int_CAND3_TLSTR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I7_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx42928z2),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p0_int[24]),.T1I1(lint_WDATA_int[24]),.T1I2(nx34006z2),.T1I3(GND),.TB1S(GND),.Q1Z(m0_oper0_wdata_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_I7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[29]),.Q1EN(tcdm_valid_p0_int_CAND3_TLSTR_9_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_9_padClk),.QRT(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[28]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[26]),.Q2EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_127_CAND4_TLSBR_9_tpGCLKBUF),.B0I1(m0_m0_control[24]),.B0I2(tcdm_result_p0[24]),.B0I3(NET_129),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.B0Z(NET_629),.Q0Z(m0_m0_control[24]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I10_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_127_CAND4_TLSBR_9_tpGCLKBUF),.T1I1(tcdm_result_p0[29]),.T1I2(NET_129),.T1I3(m0_m0_control[29]),.C1Z(NET_733),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_I10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.Q2Z(m0_m0_control[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I10_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_127_CAND4_TLSBR_9_tpGCLKBUF),.T3I1(m0_m0_control[28]),.T3I2(NET_129),.T3I3(tcdm_result_p0[28]),.C3Z(NET_710),.Q3Z(m0_m0_control[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_I11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_124),.B0I1(NET_130),.B0I2(m0_m0_dataout_int[24]),.B0I3(m1_ram_control[24]),.CD0S(VCC),.Q0DI(lint_WDATA_int[26]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.B0Z(NET_627),.Q0Z(m0_m0_control[26]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I11_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_629),.T1I1(NET_628),.T1I2(NET_627),.T1I3(NET_630),.C1Z(NET_617),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_I11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper0_wdsel_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I11_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[24]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p0[26]),.T3I1(NET_129),.T3I2(NET_127_CAND4_TLSBR_9_tpGCLKBUF),.T3I3(m0_m0_control[26]),.C3Z(NET_668),.Q3Z(m1_ram_control[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_I12_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(m1_oper0_wdsel_dup_0),.B0I1(NET_131),.B0I2(m1_m1_mode_dup_0[0]),.B0I3(NET_130),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(GND),.T0I0(NET_317),.T0I1(NET_320),.T0I2(NET_319),.T0I3(NET_318),.TB0S(GND),.B0Z(NET_320),.C0Z(NET_306),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_REQ_int),.Q2EN(RESET_int[0]),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(GND),.Q2Z(saved_REQ),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I12_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(GND),.QST(GND),.T3I0(NET_124),.T3I1(m0_m0_dataout_int[12]),.T3I2(NET_125),.T3I3(m1_m0_dataout_int[12]),.C3Z(NET_318),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_I13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001000000000000),.B0I0(GND),.B0I1(GND),.B0I2(NET_87),.B0I3(lint_BE_int[1]),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.B0Z(nx58361z1),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx19381z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_control[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx12574z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.Q2Z(m0_m0_outsel_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I13_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[13]),.Q3EN(nx58361z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_124),.T3I1(NET_125),.T3I2(m0_m0_dataout_int[17]),.T3I3(m1_m0_dataout_int[17]),.TB3S(GND),.C3Z(NET_444),.Q3Z(m0_m0_mode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_I14_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000010000000000),.B0I0(GND),.B0I1(lint_BE_int[0]),.B0I2(GND),.B0I3(NET_87),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx32122z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T0I0(NET_604),.T0I1(NET_603),.T0I2(NET_606),.T0I3(NET_605),.TB0S(GND),.B0Z(nx12574z1),.C0Z(NET_592),.Q0Z(m1_m1_control[19]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx12574z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.Q1Z(m0_m0_outsel_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I14_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000001000),.B2I0(NET_80),.B2I1(lint_BE_int[0]),.B2I2(GND),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(NET_131),.T2I1(m1_m0_control[19]),.T2I2(NET_128),.T2I3(m1_m1_control[19]),.TB2S(GND),.B2Z(nx36875z1),.C2Z(NET_491),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx12574z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_outsel_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I15_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T0I0(NET_491),.T0I1(NET_492),.T0I2(NET_494),.T0I3(NET_493),.TB0S(GND),.C0Z(NET_488),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I15_1 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx41096z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_29),.T1I1(lint_ADDR_int[11]),.T1I2(NET_34),.T1I3(GND),.C1Z(NET_130),.Q1Z(m1_m1_control[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_I15_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_131),.B2I1(m1_oper1_wmode_dup_0[1]),.B2I2(NET_130),.B2I3(m1_m1_control[7]),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[79]),.T2I1(m0_m0_dataout_int[15]),.T2I2(NET_36),.T2I3(NET_41),.TB2S(GND),.B2Z(NET_606),.C2Z(NET_402),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I15_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_130),.T3I1(NET_131),.T3I2(m1_oper1_wmode_dup_0[0]),.T3I3(m1_m1_tc_dup_0),.C3Z(NET_806),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_I16_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T0I0(m0_m0_dataout_int[13]),.T0I1(NET_41),.T0I2(fpgaio_in_int[77]),.T0I3(NET_36),.TB0S(GND),.C0Z(NET_334),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I16_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx41096z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_371),.T1I1(NET_370),.T1I2(NET_373),.T1I3(NET_372),.TB1S(GND),.C1Z(NET_353),.Q1Z(m1_m1_control[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_I16_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_m1_control[5]),.B2I1(NET_37),.B2I2(fpgaio_in_int[69]),.B2I3(NET_36),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx41096z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[65]),.T2I1(NET_37),.T2I2(m1_m1_control[1]),.T2I3(NET_36),.TB2S(GND),.B2Z(NET_828),.C2Z(NET_15),.Q2Z(m1_m1_control[5]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_I16_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx41096z1),.QCK(CLK_int_0__CAND0_TLSBR_9_padClk),.QRT(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_dataout_int[14]),.T3I1(NET_41),.T3I2(NET_36),.T3I3(fpgaio_in_int[78]),.TB3S(GND),.C3Z(NET_373),.Q3Z(m1_m1_tc_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_I17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_18),.B0I1(NET_17),.B0I2(NET_15),.B0I3(NET_16),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B0Z(NET_12),.Q0Z(m1_m1_control[30]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_757),.B1I1(NET_754),.B1I2(NET_756),.B1I3(NET_755),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(NET_756),.T1I1(NET_755),.T1I2(NET_757),.T1I3(NET_754),.TB1S(NET_758),.C1Z(NET_749),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_I17_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_37),.B2I1(m1_m1_control[30]),.B2I2(NET_66),.B2I3(m1_m0_dataout_int[30]),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T2I0(NET_37),.T2I1(NET_66),.T2I2(m1_m0_dataout_int[27]),.T2I3(m1_m1_control[27]),.TB2S(GND),.B2Z(NET_757),.C2Z(NET_685),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_control[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[7]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[71]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[69]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[75]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q3Z(fpgaio_out_dup_0[66]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q1Z(fpgaio_out_dup_0[79]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_142),.B0I1(fpgaio_in_int[58]),.B0I2(NET_114),.B0I3(m0_ram_control[26]),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B0Z(NET_659),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q3Z(m0_ram_control[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx58361z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q0Z(m0_m0_osel_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx58361z1),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_csel_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I22_0 (.tFragBitInfo(16'b0101000101000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(nx22245z2),.T0I2(lint_WDATA_int[1]),.T0I3(tcdm_rdata_p2_int[1]),.TB0S(GND),.Q0Z(m1_oper0_wdata_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I23_0 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p2_int[16]),.T0I1(GND),.T0I2(nx22245z2),.T0I3(lint_WDATA_int[16]),.TB0S(GND),.Q0Z(m1_oper0_wdata_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I24_1 (.tFragBitInfo(16'b0011001000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T1I0(nx22245z2),.T1I1(GND),.T1I2(tcdm_rdata_p2_int[26]),.T1I3(lint_WDATA_int[26]),.TB1S(GND),.Q1Z(m1_oper0_wdata_dup_0[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_I24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_I24_3 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSTR_9_padClk),.QRT(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF),.QST(GND),.T3I0(nx22245z2),.T3I1(tcdm_rdata_p2_int[4]),.T3I2(lint_WDATA_int[4]),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper0_wdata_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_I25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I25_2 (.tFragBitInfo(16'b0101000001000100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx12783z2),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(tcdm_rdata_p2_int[29]),.T2I2(lint_WDATA_int[29]),.T2I3(nx22245z2),.TB2S(GND),.Q2Z(m1_oper0_wdata_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_I25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_I26_0 (.tFragBitInfo(16'b0010001011110000),.bFragBitInfo(16'b1100010011110101),.B0I0(p2_fsm[4]),.B0I1(launch_p2),.B0I2(tcdm_valid_p2_int),.B0I3(p2_fsm[0]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx39673z1),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.T0I0(NET_165),.T0I1(NET_164),.T0I2(p2_fsm[3]),.T0I3(p2_fsm[2]),.TB0S(GND),.B0Z(NET_549),.C0Z(nx43661z1),.Q0Z(p2_fsm[4]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I26_1 (.tFragBitInfo(16'b0001000100010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.T1I0(tcdm_gnt_p2_int),.T1I1(GND),.T1I2(p2_fsm[3]),.T1I3(p2_fsm[2]),.TB1S(GND),.C1Z(NET_231),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_I26_2 (.tFragBitInfo(16'b0000010011001100),.bFragBitInfo(16'b0000110011001100),.B2I0(NET_165),.B2I1(NET_549),.B2I2(p2_fsm[3]),.B2I3(NET_231),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(NET_165),.T2I1(NET_549),.T2I2(p2_fsm[3]),.T2I3(NET_231),.TB2S(NET_164),.C2Z(nx39673z1),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I26_3 (.tFragBitInfo(16'b0000000000000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(p2_fsm[4]),.T3I1(RESET_int[0]),.T3I2(NET_231),.T3I3(p2_fsm[1]),.TB3S(GND),.C3Z(NET_230),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_I27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_I27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_I27_2 (.tFragBitInfo(16'b0000000000001100),.bFragBitInfo(16'b1111111101000000),.B2I0(NET_164),.B2I1(p2_fsm[4]),.B2I2(NET_165),.B2I3(p2_fsm[0]),.CD2S(GND),.Q2EN(nx39673z1),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(nx42664z1),.T2I2(GND),.T2I3(not_tcdm_wen_p2),.TB2S(GND),.B2Z(nx42664z1),.Q2Z(p2_fsm[3]),.B2CO(),.C2Z(),.Q2DI(GND),.T2CO());

	LOGIC_3 QL_INST_I27_3 (.tFragBitInfo(16'b0111001100000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF),.QST(GND),.T3I0(NET_164),.T3I1(p2_fsm[2]),.T3I2(NET_165),.T3I3(NET_230),.C3Z(nx20942z2),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_I28_0 (.tFragBitInfo(16'b0000011000001010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(GND),.QST(GND),.T0I0(p2_cnt[11]),.T0I1(NET_255),.T0I2(p2_fsm[0]),.T0I3(p2_cnt[10]),.TB0S(GND),.Q0Z(p2_cnt[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_I28_1 (.tFragBitInfo(16'b0000000100000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(GND),.QST(GND),.T1I0(NET_255),.T1I1(GND),.T1I2(p2_fsm[0]),.T1I3(p2_cnt[10]),.TB1S(GND),.Q1Z(p2_cnt[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_I28_2 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0000000000000001),.B2I0(p2_cnt[11]),.B2I1(p2_cnt[8]),.B2I2(p2_cnt[9]),.B2I3(p2_cnt[10]),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(GND),.QST(GND),.T2I0(GND),.T2I1(NET_208),.T2I2(p2_cnt[8]),.T2I3(p2_cnt[9]),.TB2S(GND),.B2Z(NET_165),.C2Z(NET_255),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_I28_3 (.tFragBitInfo(16'b0000011100001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx20942z2),.QCK(CLK_int_0__CAND0_BLSBR_9_padClk),.QRT(GND),.QST(GND),.T3I0(p2_cnt[8]),.T3I1(NET_208),.T3I2(p2_fsm[0]),.T3I3(p2_cnt[9]),.TB3S(GND),.Q3Z(p2_cnt[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_J3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J3_2 (.tFragBitInfo(16'b0001000100010000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2EN(nx18527z1),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.T2I0(GND),.T2I1(GND),.T2I2(nx11313z5),.T2I3(nx18527z8),.TB2S(GND),.Q2Z(p0_fsm[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.Q2DI(GND),.T2CO());

	LOGIC_3 QL_INST_J3_3 (.tFragBitInfo(16'b0000000011010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.T3I0(NET_188),.T3I1(NET_187),.T3I2(p0_fsm[4]),.T3I3(GND),.C3Z(nx18527z8),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J4_0 (.tFragBitInfo(16'b0000000000001010),.bFragBitInfo(16'b0001000000110011),.B0I0(NET_187),.B0I1(p0_fsm[1]),.B0I2(NET_188),.B0I3(p0_fsm[2]),.CD0S(GND),.Q0EN(nx18527z1),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.T0I0(p0_fsm[0]),.T0I1(GND),.T0I2(GND),.T0I3(tcdm_wen_p0_dup_0),.TB0S(GND),.B0Z(NET_186),.Q0Z(p0_fsm[1]),.B0CO(),.C0Z(),.Q0DI(GND),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J4_1 (.tFragBitInfo(16'b0000000000001110),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1EN(nx18527z1),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.T1I0(nx20521z1),.T1I1(p0_fsm[1]),.T1I2(GND),.T1I3(GND),.TB1S(GND),.Q1Z(p0_fsm[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.Q1DI(GND),.T1CO());

	LOGIC_2 QL_INST_J4_2 (.tFragBitInfo(16'b0001000100010000),.bFragBitInfo(16'b0010001100000000),.B2I0(NET_187),.B2I1(GND),.B2I2(NET_188),.B2I3(p0_fsm[2]),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.T2I0(tcdm_gnt_p0_int),.T2I1(GND),.T2I2(p0_fsm[2]),.T2I3(p0_fsm[3]),.TB2S(GND),.B2Z(nx11313z5),.C2Z(NET_217),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J4_3 (.tFragBitInfo(16'b0100111101000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx18527z1),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_187),.T3I1(NET_188),.T3I2(p0_fsm[2]),.T3I3(p0_fsm[3]),.TB3S(GND),.C3Z(nx22515z1),.Q3Z(p0_fsm[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_J6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_69),.B0I1(fpgaio_in_int[25]),.B0I2(m0_m1_dataout_int[25]),.B0I3(NET_242),.B0Z(NET_640),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J6_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_69),.T3I1(fpgaio_in_int[27]),.T3I2(m0_m1_dataout_int[27]),.T3I3(NET_242),.C3Z(NET_682),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[18]),.Q0EN(tcdm_valid_p0_int_CAND3_TLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J7_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_69),.T1I1(m0_m1_dataout_int[30]),.T1I2(NET_242),.T1I3(fpgaio_in_int[30]),.C1Z(NET_754),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[7]),.Q2EN(tcdm_valid_p0_int_CAND3_TLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[6]),.Q1EN(tcdm_valid_p0_int_CAND3_TLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_10_padClk),.QRT(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(m0_m1_tc_dup_0),.B0I1(NET_127_CAND4_TLSBR_10_tpGCLKBUF),.B0I2(NET_126_CAND3_TLSBR_10_tpGCLKBUF),.B0I3(tcdm_result_p0[6]),.B0Z(NET_805),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J10_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(tcdm_result_p0[7]),.T3I1(NET_127_CAND4_TLSBR_10_tpGCLKBUF),.T3I2(NET_126_CAND3_TLSBR_10_tpGCLKBUF),.T3I3(m0_m1_control[7]),.TB3S(GND),.C3Z(NET_605),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_J11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[17]),.Q0EN(nx49703z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.Q0Z(m0_m1_clr_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J11_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_126_CAND3_TLSBR_10_tpGCLKBUF),.T1I1(m1_m0_control[29]),.T1I2(m0_m1_control[29]),.T1I3(NET_128),.C1Z(NET_732),.Q1Z(m0_m1_control[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[29]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_control[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J11_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_126_CAND3_TLSBR_10_tpGCLKBUF),.T3I1(NET_130),.T3I2(m1_ram_control[17]),.T3I3(m0_m1_clr_dup_0),.TB3S(GND),.C3Z(NET_446),.Q3Z(m1_ram_control[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_J12_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(tcdm_result_p2[18]),.B0I1(tcdm_result_p0[18]),.B0I2(NET_127_CAND4_TLSBR_10_tpGCLKBUF),.B0I3(NET_106),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T0I0(NET_475),.T0I1(NET_476),.T0I2(NET_477),.T0I3(NET_474),.TB0S(GND),.B0Z(NET_476),.C0Z(NET_478),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J12_1 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[28]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(NET_80),.T1I2(GND),.T1I3(lint_BE_int[3]),.C1Z(nx28356z1),.Q1Z(m1_m0_control[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m0_m1_control[28]),.B2I1(NET_128),.B2I2(NET_126_CAND3_TLSBR_10_tpGCLKBUF),.B2I3(m1_m0_control[28]),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.B2Z(NET_709),.Q2Z(m0_m1_control[28]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[16]),.Q3EN(nx19381z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.Q3Z(m1_m0_rnd_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B0I0(NET_71),.B0I1(lint_ADDR_int[11]),.B0I2(GND),.B0I3(NET_33_CAND2_TLSBR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.B0Z(NET_128),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J13_1 (.tFragBitInfo(16'b0101111111111111),.bFragBitInfo(16'b0011001101111111),.B1I0(m1_m0_control[20]),.B1I1(NET_33_CAND2_TLSBR_10_tpGCLKBUF),.B1I2(NET_71),.B1I3(NET_30_CAND5_TLSBR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_71),.T1I1(NET_30_CAND5_TLSBR_10_tpGCLKBUF),.T1I2(m1_m0_control[20]),.T1I3(NET_33_CAND2_TLSBR_10_tpGCLKBUF),.TB1S(fpgaio_in_int[20]),.C1Z(NET_518),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_J13_2 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'b0000000000001000),.B2I0(lint_BE_int[2]),.B2I1(NET_87),.B2I2(GND),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_BE_int[2]),.T2I2(NET_80),.T2I3(GND),.TB2S(GND),.B2Z(nx1800z1),.C2Z(nx19381z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J13_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[20]),.Q3EN(nx19381z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_446),.T3I1(NET_444),.T3I2(NET_443),.T3I3(NET_445),.C3Z(NET_440),.Q3Z(m1_m0_control[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_804),.B0I1(NET_805),.B0I2(NET_803),.B0I3(NET_806),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.B0Z(NET_792),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J14_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T1I0(m0_m0_dataout_int[7]),.T1I1(m1_m0_dataout_int[7]),.T1I2(NET_124),.T1I3(NET_125),.C1Z(NET_604),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J14_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_125),.B2I1(m1_m0_dataout_int[6]),.B2I2(NET_124),.B2I3(m0_m0_dataout_int[6]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T2I0(NET_489),.T2I1(NET_488),.T2I2(NET_486),.T2I3(NET_487),.TB2S(GND),.B2Z(NET_804),.Q2Z(lint_RDATA_dup_0[19]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_J14_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T3I0(NET_439),.T3I1(NET_438),.T3I2(NET_440),.T3I3(NET_441),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_J15_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000100000000),.B0I0(GND),.B0I1(GND),.B0I2(lint_ADDR_int[9]),.B0I3(NET_82),.CD0S(VCC),.Q0DI(lint_WDATA_int[19]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T0I0(NET_126_CAND3_TLSBR_10_tpGCLKBUF),.T0I1(NET_130),.T0I2(m0_m1_sat_dup_0),.T0I3(m1_ram_control[18]),.TB0S(GND),.B0Z(NET_570),.C0Z(NET_474),.Q0Z(m1_ram_control[19]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J15_1 (.tFragBitInfo(16'b0111111101111111),.bFragBitInfo(16'b0001001111111111),.B1I0(NET_71),.B1I1(NET_30_CAND5_TLSBR_10_tpGCLKBUF),.B1I2(m1_m0_outsel_dup_0[1]),.B1I3(NET_33_CAND2_TLSBR_10_tpGCLKBUF),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(m1_m0_outsel_dup_0[1]),.T1I1(NET_33_CAND2_TLSBR_10_tpGCLKBUF),.T1I2(NET_71),.T1I3(NET_30_CAND5_TLSBR_10_tpGCLKBUF),.TB1S(fpgaio_in_int[1]),.C1Z(NET_68),.Q1Z(m1_ram_control[18]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_J15_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000010000000000),.B2I0(GND),.B2I1(NET_33_CAND2_TLSBR_10_tpGCLKBUF),.B2I2(GND),.B2I3(NET_30_CAND5_TLSBR_10_tpGCLKBUF),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx49703z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T2I0(NET_126_CAND3_TLSBR_10_tpGCLKBUF),.T2I1(m1_ram_control[19]),.T2I2(m0_m1_control[19]),.T2I3(NET_130),.TB2S(GND),.B2Z(NET_242),.C2Z(NET_494),.Q2Z(m0_m1_control[19]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_J15_3 (.tFragBitInfo(16'b0111111101111111),.bFragBitInfo(16'b0001001111111111),.B3I0(NET_71),.B3I1(NET_30_CAND5_TLSBR_10_tpGCLKBUF),.B3I2(m1_m0_outsel_dup_0[4]),.B3I3(NET_33_CAND2_TLSBR_10_tpGCLKBUF),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx49703z1),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_outsel_dup_0[4]),.T3I1(NET_33_CAND2_TLSBR_10_tpGCLKBUF),.T3I2(NET_71),.T3I3(NET_30_CAND5_TLSBR_10_tpGCLKBUF),.TB3S(fpgaio_in_int[4]),.C3Z(NET_867),.Q3Z(m0_m1_sat_dup_0),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_J16_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_825),.B0I1(NET_826),.B0I2(NET_824),.B0I3(NET_823),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T0I0(NET_825),.T0I1(NET_826),.T0I2(NET_824),.T0I3(NET_823),.TB0S(NET_827),.Q0Z(lint_RDATA_dup_0[5]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_684),.B1I1(NET_683),.B1I2(NET_685),.B1I3(NET_682),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T1I0(NET_685),.T1I1(NET_682),.T1I2(NET_684),.T1I3(NET_683),.TB1S(NET_686),.C1Z(NET_677),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_J16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000001000000),.B2I0(lint_ADDR_int[3]),.B2I1(lint_ADDR_int[5]),.B2I2(lint_ADDR_int[6]),.B2I3(lint_ADDR_int[4]),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.B2Z(NET_30),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J16_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF),.T3I0(NET_36),.T3I1(m0_m0_dataout_int[4]),.T3I2(fpgaio_in_int[68]),.T3I3(NET_41),.C3Z(NET_852),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_643),.B0I1(NET_641),.B0I2(NET_640),.B0I3(NET_642),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[18]),.Q0EN(tcdm_valid_p2_int_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T0I0(NET_643),.T0I1(NET_641),.T0I2(NET_640),.T0I3(NET_642),.TB0S(NET_644),.C0Z(NET_635),.Q0Z(tcdm_result_p2[18]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J17_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_37),.T1I1(m1_m0_dataout_int[25]),.T1I2(NET_66),.T1I3(m1_m1_control[25]),.C1Z(NET_643),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_J17_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B2I0(fpgaio_in_int[73]),.B2I1(NET_36),.B2I2(m0_m0_dataout_int[9]),.B2I3(NET_41),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_in_int[72]),.T2I1(NET_36),.T2I2(NET_41),.T2I3(m0_m0_dataout_int[8]),.TB2S(GND),.B2Z(NET_235),.C2Z(NET_381),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_J17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[25]),.Q3EN(nx23147z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_control[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_144),.B0I1(fpgaio_in_int[24]),.B0I2(NET_143),.B0I3(m1_m1_dataout_int[24]),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B0Z(NET_621),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010101000000000),.B1I0(NET_724),.B1I1(tcdm_result_p2[29]),.B1I2(NET_106),.B1I3(NET_723),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_106),.T1I1(NET_723),.T1I2(NET_724),.T1I3(tcdm_result_p2[29]),.TB1S(NET_725),.C1Z(NET_720),.Q1Z(fpgaio_out_dup_0[67]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_J18_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_144),.B2I1(m1_m1_dataout_int[29]),.B2I2(fpgaio_in_int[29]),.B2I3(NET_143),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T2I0(NET_144),.T2I1(m1_m1_dataout_int[26]),.T2I2(NET_143),.T2I3(fpgaio_in_int[26]),.TB2S(GND),.B2Z(NET_725),.C2Z(NET_660),.Q2Z(fpgaio_out_dup_0[68]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_J18_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_144),.T3I1(fpgaio_in_int[28]),.T3I2(NET_143),.T3I3(m1_m1_dataout_int[28]),.C3Z(NET_702),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000011000000),.B1I0(tcdm_result_p2[24]),.B1I1(NET_619),.B1I2(NET_620),.B1I3(NET_106),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T1I0(NET_620),.T1I1(NET_106),.T1I2(tcdm_result_p2[24]),.T1I3(NET_619),.TB1S(NET_621),.C1Z(NET_616),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_J19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010101000000000),.B2I0(NET_659),.B2I1(tcdm_result_p2[26]),.B2I2(NET_106),.B2I3(NET_658),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T2I0(NET_659),.T2I1(tcdm_result_p2[26]),.T2I2(NET_106),.T2I3(NET_658),.TB2S(NET_660),.C2Z(NET_655),.Q2Z(fpgaio_out_dup_0[78]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_J19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010101000000000),.B3I0(NET_700),.B3I1(tcdm_result_p2[28]),.B3I2(NET_106),.B3I3(NET_701),.CD3S(VCC),.Q3DI(lint_WDATA_int[6]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_106),.T3I1(NET_701),.T3I2(NET_700),.T3I3(tcdm_result_p2[28]),.TB3S(NET_702),.C3Z(NET_697),.Q3Z(m1_oper1_wmode_dup_0[0]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_J20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[28]),.Q0EN(tcdm_valid_p2_int_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p2[28]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J20_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_28),.T3I1(m0_m0_outsel_dup_0[3]),.T3I2(fpgaio_in_int[35]),.T3I3(NET_27_CAND5_BLSTR_10_tpGCLKBUF),.C3Z(NET_875),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_J21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_J21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[24]),.Q1EN(tcdm_valid_p2_int_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[26]),.Q2EN(tcdm_valid_p2_int_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p2[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J22_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T0I0(NET_79),.T0I1(NET_6),.T0I2(NET_8),.T0I3(lint_ADDR_int[14]),.TB0S(GND),.C0Z(NET_482),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J22_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[29]),.Q1EN(tcdm_valid_p2_int_CAND2_BLSTR_10_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[14]),.T1I1(NET_6),.T1I2(NET_8),.T1I3(NET_10),.TB1S(GND),.C1Z(nx22245z2),.Q1Z(tcdm_result_p2[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_J22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_J22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[3]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_10_padClk),.QRT(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF),.QST(GND),.Q3Z(m1_oper0_wmode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_J26_0 (.tFragBitInfo(16'b0000000000001110),.bFragBitInfo(16'b0000000000000001),.B0I0(p2_fsm[1]),.B0I1(GND),.B0I2(GND),.B0I3(p2_fsm[0]),.CD0S(GND),.Q0EN(nx39673z1),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T0I0(p2_fsm[1]),.T0I1(nx41667z1),.T0I2(GND),.T0I3(GND),.TB0S(GND),.B0Z(NET_163),.Q0Z(p2_fsm[2]),.B0CO(),.C0Z(),.Q0DI(GND),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J26_1 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(tcdm_valid_p2_int),.T1I2(p2_fsm[4]),.T1I3(tcdm_wen_p2_dup_0),.TB1S(GND),.C1Z(nx22245z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_J26_2 (.tFragBitInfo(16'b0000000001010000),.bFragBitInfo(16'b0000000000100000),.B2I0(NET_165),.B2I1(NET_164),.B2I2(p2_fsm[4]),.B2I3(tcdm_wen_p2_dup_0),.CD2S(GND),.Q2EN(nx39673z1),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(GND),.T2I2(p2_fsm[0]),.T2I3(tcdm_wen_p2_dup_0),.TB2S(GND),.B2Z(nx41667z1),.Q2Z(p2_fsm[1]),.B2CO(),.C2Z(),.Q2DI(GND),.T2CO());

	LOGIC_3 QL_INST_J26_3 (.tFragBitInfo(16'b0101010111110101),.bFragBitInfo(16'b0010111110101111),.B3I0(NET_163),.B3I1(p2_fsm[2]),.B3I2(NET_162),.B3I3(NET_164),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.QST(GND),.T3I0(NET_162),.T3I1(NET_164),.T3I2(NET_163),.T3I3(p2_fsm[2]),.TB3S(NET_165),.C3Z(nx11311z2),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_J27_0 (.tFragBitInfo(16'b0010000000100010),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.T0I0(p2_fsm[4]),.T0I1(GND),.T0I2(NET_164),.T0I3(NET_165),.TB0S(GND),.C0Z(nx39673z6),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_J27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_J27_2 (.tFragBitInfo(16'b0000001100000010),.bFragBitInfo(16'b0010000000100010),.B2I0(p2_fsm[2]),.B2I1(GND),.B2I2(NET_164),.B2I3(NET_165),.CD2S(GND),.Q2EN(nx39673z1),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.T2I0(nx11311z3),.T2I1(GND),.T2I2(GND),.T2I3(nx39673z6),.TB2S(GND),.B2Z(nx11311z3),.Q2Z(p2_fsm[0]),.B2CO(),.C2Z(),.Q2DI(GND),.T2CO());

	LOGIC_3 QL_INST_J27_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_10_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF),.T3I0(tcdm_wen_p2_dup_0),.T3I1(GND),.T3I2(GND),.T3I3(GND),.C3Z(not_tcdm_wen_p2),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_K4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[26]),.Q1EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[28]),.Q3EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[29]),.Q1EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[21]),.Q1EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_11_padClk),.QRT(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[31]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx57183z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_tc_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx57183z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_control[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.Q0Z(m1_m0_control[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[24]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_control[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_128),.B2I1(m1_m0_control[26]),.B2I2(m0_m1_control[26]),.B2I3(NET_126_CAND3_TLSBR_11_tpGCLKBUF),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx28356z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.B2Z(NET_667),.Q2Z(m1_m0_control[26]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K11_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[26]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(NET_128),.T3I1(m1_m0_control[24]),.T3I2(m0_m1_control[24]),.T3I3(NET_126_CAND3_TLSBR_11_tpGCLKBUF),.C3Z(NET_628),.Q3Z(m0_m1_control[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_K12_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_32),.B0I1(NET_571),.B0I2(lint_BE_int[0]),.B0I3(NET_257),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(m1_m0_mode_dup_0[0]),.T0I1(NET_128),.T0I2(NET_129),.T0I3(m0_m0_mode_dup_0[0]),.TB0S(GND),.B0Z(nx57183z1),.C0Z(NET_317),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx23147z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_reset_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K12_2 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b1000000000000000),.B2I0(lint_BE_int[3]),.B2I1(NET_571),.B2I2(NET_257),.B2I3(NET_32),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_80),.T2I1(lint_BE_int[1]),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(nx40728z1),.C2Z(nx10406z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K12_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(NET_32),.T3I1(NET_571),.T3I2(lint_BE_int[2]),.T3I3(NET_257),.C3Z(nx49703z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_K13_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0001000000000000),.B0I0(GND),.B0I1(GND),.B0I2(NET_87),.B0I3(lint_BE_int[3]),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(NET_32),.T0I1(NET_257),.T0I2(NET_258),.T0I3(lint_BE_int[3]),.TB0S(GND),.B0Z(nx10775z1),.C0Z(nx23147z1),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K13_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_257),.T1I1(NET_32),.T1I2(NET_258),.T1I3(lint_BE_int[2]),.C1Z(nx32122z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_257),.B2I1(lint_BE_int[1]),.B2I2(NET_258),.B2I3(NET_32),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.B2Z(nx41097z1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K13_3 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0000011111111111),.B3I0(fpgaio_in_int[31]),.B3I1(NET_30_CAND5_TLSBR_11_tpGCLKBUF),.B3I2(saved_REQ),.B3I3(NET_33_CAND2_TLSBR_11_tpGCLKBUF),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx58361z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(saved_REQ),.T3I1(NET_33_CAND2_TLSBR_11_tpGCLKBUF),.T3I2(fpgaio_in_int[31]),.T3I3(NET_30_CAND5_TLSBR_11_tpGCLKBUF),.TB3S(NET_40),.C3Z(NET_924),.Q3Z(m0_m0_mode_dup_0[0]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_82),.B0I1(NET_32),.B0I2(NET_83),.B0I3(NET_81),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx41097z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T0I0(NET_82),.T0I1(NET_32),.T0I2(NET_83),.T0I3(NET_81),.TB0S(NET_31),.C0Z(NET_87),.Q0Z(m1_m1_control[11]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K14_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_124),.T1I1(m0_m0_dataout_int[2]),.T1I2(m1_m0_dataout_int[2]),.T1I3(NET_125),.C1Z(NET_906),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K14_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000001000000),.B2I0(GND),.B2I1(NET_38),.B2I2(lint_ADDR_int[2]),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_257),.T2I1(NET_32),.T2I2(NET_258),.T2I3(lint_BE_int[0]),.TB2S(GND),.B2Z(NET_258),.C2Z(nx41096z1),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_83),.B3I1(NET_81),.B3I2(NET_82),.B3I3(NET_32),.CD3S(VCC),.Q3DI(lint_WDATA_int[12]),.Q3EN(nx10406z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(NET_82),.T3I1(NET_32),.T3I2(NET_83),.T3I3(NET_81),.TB3S(NET_38),.C3Z(NET_80),.Q3Z(m1_m0_mode_dup_0[0]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(m0_m0_dataout_int[0]),.B0I1(NET_125),.B0I2(m1_m0_dataout_int[0]),.B0I3(NET_124),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.B0Z(NET_121),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K15_1 (.tFragBitInfo(16'b0111011111111111),.bFragBitInfo(16'b0001010111111111),.B1I0(m1_m0_mode_dup_0[1]),.B1I1(fpgaio_in_int[13]),.B1I2(NET_30_CAND5_TLSBR_11_tpGCLKBUF),.B1I3(NET_33_CAND2_TLSBR_11_tpGCLKBUF),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx10406z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_30_CAND5_TLSBR_11_tpGCLKBUF),.T1I1(NET_33_CAND2_TLSBR_11_tpGCLKBUF),.T1I2(m1_m0_mode_dup_0[1]),.T1I3(fpgaio_in_int[13]),.TB1S(NET_71),.C1Z(NET_917),.Q1Z(m1_m0_mode_dup_0[1]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_K15_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_35),.B2I1(NET_39),.B2I2(lint_ADDR_int[11]),.B2I3(NET_38),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_35),.T2I1(NET_39),.T2I2(GND),.T2I3(NET_38),.TB2S(GND),.B2Z(NET_131),.C2Z(NET_37),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K15_3 (.tFragBitInfo(16'b0111011111111111),.bFragBitInfo(16'b0001111101011111),.B3I0(m1_m0_control[9]),.B3I1(NET_30_CAND5_TLSBR_11_tpGCLKBUF),.B3I2(NET_33_CAND2_TLSBR_11_tpGCLKBUF),.B3I3(fpgaio_in_int[9]),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx10406z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(NET_33_CAND2_TLSBR_11_tpGCLKBUF),.T3I1(fpgaio_in_int[9]),.T3I2(m1_m0_control[9]),.T3I3(NET_30_CAND5_TLSBR_11_tpGCLKBUF),.TB3S(NET_71),.C3Z(NET_914),.Q3Z(m1_m0_control[9]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B0I0(NET_29),.B0I1(GND),.B0I2(GND),.B0I3(NET_30_CAND5_TLSBR_11_tpGCLKBUF),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx58361z1),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.B0Z(NET_28),.Q0Z(m0_m0_control[11]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K16_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T1I0(NET_33_CAND2_TLSBR_11_tpGCLKBUF),.T1I1(GND),.T1I2(NET_38),.T1I3(NET_57),.TB1S(GND),.C1Z(NET_55),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_K16_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_829),.B2I1(NET_828),.B2I2(NET_830),.B2I3(NET_831),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T2I0(m0_m0_control[11]),.T2I1(NET_27),.T2I2(NET_37),.T2I3(m1_m1_control[11]),.TB2S(GND),.B2Z(NET_824),.C2Z(NET_292),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_K16_3 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_11_padClk),.QRT(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[4]),.T3I1(GND),.T3I2(lint_ADDR_int[3]),.T3I3(GND),.TB3S(GND),.C3Z(NET_38),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_K17_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B0I0(NET_284),.B0I1(NET_282),.B0I2(NET_283),.B0I3(NET_281),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z66),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.T0I0(NET_284),.T0I1(NET_282),.T0I2(NET_283),.T0I3(NET_281),.TB0S(NET_285),.Q0Z(lint_RDATA_dup_0[11]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K17_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.T1I0(NET_292),.T1I1(NET_930),.T1I2(NET_294),.T1I3(NET_295),.C1Z(NET_283),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_K17_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z66),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.T2I0(NET_259),.T2I1(NET_262),.T2I2(NET_260),.T2I3(NET_261),.TB2S(GND),.Q2Z(lint_RDATA_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_K17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q0Z(fpgaio_out_dup_0[73]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K18_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[6]),.Q1EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_in_int[43]),.T1I1(fpgaio_in_int[11]),.T1I2(NET_28),.T1I3(NET_242),.TB1S(GND),.C1Z(NET_296),.Q1Z(fpgaio_out_dup_0[70]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_K18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[72]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K18_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[4]),.T3I1(NET_204),.T3I2(lint_ADDR_int[6]),.T3I3(NET_93),.C3Z(nx58292z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_K19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx53524z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q2Z(fpgaio_out_dup_0[76]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K19_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[6]),.T3I1(NET_204),.T3I2(NET_93),.T3I3(lint_ADDR_int[4]),.C3Z(nx53524z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_K20_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0101011111011111),.B0I0(NET_34),.B0I1(lint_ADDR_int_2__CAND3_BLSTR_11_tpGCLKBUF),.B0I2(m0_coef_rmode_dup_0[1]),.B0I3(m1_coef_rmode_dup_0[1]),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx58361z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T0I0(NET_34),.T0I1(lint_ADDR_int_2__CAND3_BLSTR_11_tpGCLKBUF),.T0I2(m0_coef_rmode_dup_0[1]),.T0I3(m1_coef_rmode_dup_0[1]),.TB0S(NET_35),.C0Z(NET_238),.Q0Z(m0_m0_control[10]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx58361z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q2Z(m0_m0_control[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K20_3 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0001000000110000),.B3I0(m0_m0_control[9]),.B3I1(fpgaio_in_int[41]),.B3I2(NET_238),.B3I3(NET_27_CAND5_BLSTR_11_tpGCLKBUF),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(NET_238),.T3I1(NET_27_CAND5_BLSTR_11_tpGCLKBUF),.T3I2(m0_m0_control[9]),.T3I3(fpgaio_in_int[41]),.TB3S(NET_28),.C3Z(NET_234),.Q3Z(m1_oper1_wmode_dup_0[1]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_K21_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0011101101111111),.B0I0(lint_ADDR_int_2__CAND3_BLSTR_11_tpGCLKBUF),.B0I1(NET_34),.B0I2(m1_coef_rmode_dup_0[0]),.B0I3(m0_coef_rmode_dup_0[0]),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int_2__CAND3_BLSTR_11_tpGCLKBUF),.T0I1(NET_34),.T0I2(m1_coef_rmode_dup_0[0]),.T0I3(m0_coef_rmode_dup_0[0]),.TB0S(NET_35),.C0Z(NET_383),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_K21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[8]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_rmode_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K21_2 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0000000000101010),.B2I0(NET_833),.B2I1(NET_27_CAND5_BLSTR_11_tpGCLKBUF),.B2I2(m0_m0_outsel_dup_0[5]),.B2I3(fpgaio_in_int[37]),.CD2S(VCC),.Q2DI(lint_WDATA_int[8]),.Q2EN(nx58361z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T2I0(NET_833),.T2I1(NET_27_CAND5_BLSTR_11_tpGCLKBUF),.T2I2(m0_m0_outsel_dup_0[5]),.T2I3(fpgaio_in_int[37]),.TB2S(NET_28),.C2Z(NET_830),.Q2Z(m0_m0_control[8]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_K21_3 (.tFragBitInfo(16'b0000101010101010),.bFragBitInfo(16'b0000000001110000),.B3I0(m0_m0_control[8]),.B3I1(NET_27_CAND5_BLSTR_11_tpGCLKBUF),.B3I2(NET_383),.B3I3(fpgaio_in_int[40]),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.T3I0(NET_383),.T3I1(fpgaio_in_int[40]),.T3I2(m0_m0_control[8]),.T3I3(NET_27_CAND5_BLSTR_11_tpGCLKBUF),.TB3S(NET_28),.C3Z(NET_380),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_K22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_rmode_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_11_padClk),.QRT(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[11]),.Q0EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[29]),.Q3EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[27]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_K28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_K28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_K28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[28]),.Q2EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_K28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_11_padClk),.QRT(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[24]),.Q3EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[17]),.Q2EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[20]),.Q3EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[25]),.Q2EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_12_padClk),.QRT(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[2]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(tcdm_result_p0[2]),.B0I1(m0_m1_outsel_dup_0[2]),.B0I2(NET_126_CAND3_TLSBR_12_tpGCLKBUF),.B0I3(NET_127_CAND4_TLSBR_12_tpGCLKBUF),.B0Z(NET_907),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L11_0 (.tFragBitInfo(16'b0011111100000000),.bFragBitInfo(16'b0001010100000000),.B0I0(tcdm_result_p1[10]),.B0I1(m0_m0_dataout_int[10]),.B0I2(NET_41),.B0I3(NET_268),.T0I0(tcdm_result_p1[10]),.T0I1(m0_m0_dataout_int[10]),.T0I2(NET_41),.T0I3(NET_268),.TB0S(NET_42),.C0Z(NET_263),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_L11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m0_m0_dataout_int[5]),.B2I1(NET_42),.B2I2(NET_41),.B2I3(tcdm_result_p1[5]),.B2Z(NET_831),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L11_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(tcdm_result_p1[1]),.T3I1(m0_m0_dataout_int[1]),.T3I2(NET_41),.T3I3(NET_42),.C3Z(NET_18),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_63),.B0I1(NET_241),.B0I2(m0_m1_control[27]),.B0I3(m1_m0_control[27]),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx28356z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.B0Z(NET_678),.Q0Z(m1_m0_control[25]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L12_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_571),.T1I1(lint_BE_int[1]),.T1I2(NET_257),.T1I3(NET_32),.C1Z(nx58678z1),.Q1Z(m0_m1_control[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_L12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_control[27]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L12_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_63),.T3I1(NET_241),.T3I2(m0_m1_control[25]),.T3I3(m1_m0_control[25]),.C3Z(NET_636),.Q3Z(m1_m0_control[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L14_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[5]),.T0I1(GND),.T0I2(GND),.T0I3(lint_ADDR_int[6]),.TB0S(GND),.C0Z(NET_32),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L14_1 (.tFragBitInfo(16'b0010001000100010),.bFragBitInfo(16'b1000100011111000),.B1I0(NET_31),.B1I1(fpgaio_oe_dup_0[20]),.B1I2(NET_67),.B1I3(tcdm_be_p0_dup_0[0]),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx49703z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_67),.T1I1(tcdm_be_p0_dup_0[0]),.T1I2(NET_31),.T1I3(fpgaio_oe_dup_0[20]),.TB1S(NET_57),.C1Z(NET_920),.Q1Z(m0_m1_control[20]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_L14_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000010000000),.B2I0(NET_33_CAND2_TLSBR_12_tpGCLKBUF),.B2I1(NET_32),.B2I2(NET_31),.B2I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T2I0(m1_m0_dataout_int[20]),.T2I1(NET_66),.T2I2(NET_63),.T2I3(m0_m1_control[20]),.TB2S(GND),.B2Z(NET_129),.C2Z(NET_517),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_L14_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_32),.T3I1(NET_33_CAND2_TLSBR_12_tpGCLKBUF),.T3I2(NET_31),.T3I3(GND),.C3Z(NET_27),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L15_0 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'b0000100000000000),.B0I0(NET_31),.B0I1(NET_35),.B0I2(lint_ADDR_int[11]),.B0I3(NET_39),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T0I0(GND),.T0I1(lint_ADDR_int[6]),.T0I2(lint_ADDR_int[5]),.T0I3(lint_ADDR_int[2]),.TB0S(GND),.B0Z(NET_126),.C0Z(NET_39),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L15_1 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T1I0(NET_398),.T1I1(NET_397),.T1I2(NET_396),.T1I3(NET_395),.TB1S(GND),.Q1Z(lint_RDATA_dup_0[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_L15_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_31),.B2I1(NET_35),.B2I2(GND),.B2I3(NET_39),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T2I0(NET_402),.T2I1(NET_401),.T2I2(NET_399),.T2I3(NET_400),.TB2S(GND),.B2Z(NET_63),.C2Z(NET_396),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_L15_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.T3I0(NET_323),.T3I1(GND),.T3I2(NET_324),.T3I3(NET_322),.TB3S(GND),.C3Z(NET_307),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_L16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[27]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_ram_control[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L16_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T1I0(NET_27),.T1I1(NET_300),.T1I2(m0_m0_control[27]),.T1I3(m1_ram_control[27]),.C1Z(NET_680),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_L16_2 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_639),.B2I1(NET_638),.B2I2(NET_636),.B2I3(NET_637),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T2I0(NET_31),.T2I1(GND),.T2I2(NET_57),.T2I3(NET_29),.TB2S(GND),.B2Z(NET_634),.C2Z(NET_72),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_L16_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[27]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_12_padClk),.QRT(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF),.QST(GND),.T3I0(NET_678),.T3I1(NET_681),.T3I2(NET_680),.T3I3(NET_679),.C3Z(NET_676),.Q3Z(m0_m0_control[27]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_L17_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b1011111100111111),.B0I0(tcdm_result_p2[30]),.B0I1(NET_748),.B0I2(NET_747),.B0I3(NET_21_CAND4_BLSTR_12_tpGCLKBUF),.CD0S(GND),.Q0DI(GND),.Q0EN(nx49808z66),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.T0I0(tcdm_result_p2[30]),.T0I1(NET_748),.T0I2(NET_747),.T0I3(NET_21_CAND4_BLSTR_12_tpGCLKBUF),.TB0S(NET_749),.Q0Z(lint_RDATA_dup_0[30]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L17_1 (.tFragBitInfo(16'b1011111111111111),.bFragBitInfo(16'b0111011101111111),.B1I0(NET_40),.B1I1(NET_35),.B1I2(lint_ADDR_int_2__CAND3_BLSTR_12_tpGCLKBUF),.B1I3(fpgaio_in_int[74]),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.T1I0(lint_ADDR_int_2__CAND3_BLSTR_12_tpGCLKBUF),.T1I1(fpgaio_in_int[74]),.T1I2(NET_40),.T1I3(NET_35),.TB1S(i_events[10]),.C1Z(NET_268),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_L17_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b1101010111111111),.B2I0(NET_633),.B2I1(NET_21_CAND4_BLSTR_12_tpGCLKBUF),.B2I2(tcdm_result_p2[25]),.B2I3(NET_634),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z66),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.T2I0(NET_633),.T2I1(NET_21_CAND4_BLSTR_12_tpGCLKBUF),.T2I2(tcdm_result_p2[25]),.T2I3(NET_634),.TB2S(NET_635),.Q2Z(lint_RDATA_dup_0[25]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_L17_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b1101111101011111),.B3I0(NET_675),.B3I1(tcdm_result_p2[27]),.B3I2(NET_676),.B3I3(NET_21_CAND4_BLSTR_12_tpGCLKBUF),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z66),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.T3I0(NET_676),.T3I1(NET_21_CAND4_BLSTR_12_tpGCLKBUF),.T3I2(NET_675),.T3I3(tcdm_result_p2[27]),.TB3S(NET_677),.Q3Z(lint_RDATA_dup_0[27]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_L18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100110000000000),.B0I0(tcdm_result_p2[10]),.B0I1(NET_264),.B0I2(NET_21_CAND4_BLSTR_12_tpGCLKBUF),.B0I3(NET_263),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p2[10]),.T0I1(NET_264),.T0I2(NET_21_CAND4_BLSTR_12_tpGCLKBUF),.T0I3(NET_263),.TB0S(NET_265),.C0Z(NET_260),.Q0Z(m1_ram_control[25]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_L18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(m0_m0_control[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L18_2 (.tFragBitInfo(16'b0000011100000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_ram_control[25]),.B2I1(NET_300),.B2I2(m0_m0_control[25]),.B2I3(NET_27_CAND5_BLSTR_12_tpGCLKBUF),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[10]),.Q2EN(tcdm_valid_p2_int_CAND2_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_oe_dup_0[52]),.T2I1(NET_72),.T2I2(NET_526),.T2I3(NET_527),.TB2S(GND),.B2Z(NET_638),.C2Z(NET_521),.Q2Z(tcdm_result_p2[10]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_L18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[25]),.Q1EN(tcdm_valid_p2_int_CAND2_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[30]),.Q2EN(tcdm_valid_p2_int_CAND2_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p2[30]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[27]),.Q1EN(tcdm_valid_p2_int_CAND2_BLSTR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L20_3 (.tFragBitInfo(16'b0101000011110000),.bFragBitInfo(16'b0000000000101010),.B3I0(NET_267),.B3I1(NET_27_CAND5_BLSTR_12_tpGCLKBUF),.B3I2(m0_m0_control[10]),.B3I3(fpgaio_in_int[42]),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_control[10]),.T3I1(fpgaio_in_int[42]),.T3I2(NET_267),.T3I3(NET_27_CAND5_BLSTR_12_tpGCLKBUF),.TB3S(NET_28),.C3Z(NET_265),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_L24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx33579z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx33579z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx33579z1),.QCK(CLK_int_0__CAND0_BLSTR_12_padClk),.QRT(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[14]),.Q0EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[17]),.Q0EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[17]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[20]),.Q1EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[21]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[19]),.Q3EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[24]),.Q0EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[25]),.Q1EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L27_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_L28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_L28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_L28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[26]),.Q2EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_L28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_12_padClk),.QRT(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[10]),.Q1EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_waddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[1]),.Q3EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_waddr_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[6]),.Q0EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_waddr_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[11]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_waddr_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M4_0 (.tFragBitInfo(16'b0000000000001110),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0EN(nx11313z3),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(nx11313z1),.T0I1(nx22515z1),.T0I2(GND),.T0I3(GND),.TB0S(GND),.Q0Z(tcdm_req_p0_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.Q0DI(GND),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M4_2 (.tFragBitInfo(16'b1110111011111110),.bFragBitInfo(16'b1010101011111010),.B2I0(nx11313z1),.B2I1(NET_186),.B2I2(tcdm_gnt_p0_int),.B2I3(tcdm_fmo_p0_int),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.T2I0(nx11313z1),.T2I1(NET_186),.T2I2(tcdm_gnt_p0_int),.T2I3(tcdm_fmo_p0_int),.TB2S(p0_fsm[0]),.C2Z(nx11313z3),.Q2Z(m0_coef_wdata_dup_0[6]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_M4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_wdata_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdata_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[5]),.Q0EN(tcdm_valid_p0_int_CAND3_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wdata_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[18]),.Q3EN(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_wdata_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[15]),.Q0EN(tcdm_valid_p0_int_CAND3_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p0_int[12]),.Q2EN(tcdm_valid_p0_int_CAND3_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[14]),.Q1EN(tcdm_valid_p0_int_CAND3_TLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_13_padClk),.QRT(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[3]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_wmode_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[2]),.Q3EN(nx57183z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_outsel_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M11_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_127_CAND4_TLSBR_13_tpGCLKBUF),.T2I1(NET_126_CAND3_TLSBR_13_tpGCLKBUF),.T2I2(m0_m1_mode_dup_0[0]),.T2I3(tcdm_result_p0[12]),.TB2S(GND),.C2Z(NET_319),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_M11_3 (.tFragBitInfo(16'b0011000011110000),.bFragBitInfo(16'b0000001000001010),.B3I0(NET_878),.B3I1(NET_41),.B3I2(tcdm_result_p1[3]),.B3I3(m0_m0_dataout_int[3]),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx28356z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p1[3]),.T3I1(m0_m0_dataout_int[3]),.T3I2(NET_878),.T3I3(NET_41),.TB3S(NET_42),.C3Z(NET_876),.Q3Z(m1_m0_reset_dup_0),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_M12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.Q0Z(m0_m1_reset_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M12_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx28356z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_63),.T1I1(NET_241),.T1I2(m1_m0_reset_dup_0),.T1I3(m0_m1_reset_dup_0),.C1Z(NET_770),.Q1Z(m1_m0_control[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_M12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_63),.B2I1(NET_241),.B2I2(m1_m0_control[30]),.B2I3(m0_m1_control[30]),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B2Z(NET_750),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[30]),.Q3EN(nx40728z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_control[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_875),.B0I1(NET_876),.B0I2(NET_873),.B0I3(NET_874),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.B0Z(NET_870),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M13_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.T1I0(NET_20),.T1I1(tcdm_result_p0[3]),.T1I2(NET_293),.T1I3(m0_oper0_wmode_dup_0[1]),.C1Z(NET_873),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_M13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M13_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.T3I0(NET_869),.T3I1(NET_871),.T3I2(NET_872),.T3I3(NET_870),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_M14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1010111010101111),.B0I0(NET_783),.B0I1(NET_784),.B0I2(nx7012z2),.B0I3(NET_785),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B0Z(nx49808z66),.Q0Z(i_events[3]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M14_1 (.tFragBitInfo(16'b1101111111111111),.bFragBitInfo(16'b0011111101111111),.B1I0(fpgaio_in_int[67]),.B1I1(NET_40),.B1I2(NET_35),.B1I3(lint_ADDR_int[2]),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_35),.T1I1(lint_ADDR_int[2]),.T1I2(fpgaio_in_int[67]),.T1I3(NET_40),.TB1S(i_events[3]),.C1Z(NET_878),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_M14_2 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b0000101000001000),.B2I0(NET_82),.B2I1(NET_74),.B2I2(lint_ADDR_int[9]),.B2I3(NET_141),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_82),.T2I1(NET_83),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(NET_784),.C2Z(NET_257),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_M14_3 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_257),.T3I1(NET_1),.T3I2(GND),.T3I3(NET_141),.C3Z(nx60509z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M15_0 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'b0000000000010000),.B0I0(GND),.B0I1(GND),.B0I2(NET_86),.B0I3(lint_ADDR_int[2]),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[15]),.T0I1(GND),.T0I2(GND),.T0I3(NET_9),.TB0S(GND),.B0Z(NET_81),.C0Z(NET_6),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M15_1 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[15]),.T1I1(lint_ADDR_int[12]),.T1I2(lint_ADDR_int[14]),.T1I3(NET_9),.TB1S(GND),.C1Z(NET_211),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_M15_2 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[20]),.Q2EN(nx32122z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[15]),.T2I1(lint_ADDR_int[13]),.T2I2(lint_ADDR_int[14]),.T2I3(NET_9),.TB2S(GND),.C2Z(NET_78),.Q2Z(m1_m1_control[20]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_M15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_5),.B3I1(NET_84),.B3I2(NET_6),.B3I3(NET_83),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(NET_6),.T3I1(NET_83),.T3I2(NET_5),.T3I3(NET_84),.TB3S(NET_74),.C3Z(NET_91),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_M16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_751),.B0I1(NET_752),.B0I2(NET_753),.B0I3(NET_750),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx10775z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B0Z(NET_748),.Q0Z(m0_m0_control[30]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M16_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[30]),.Q1EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_6),.T1I1(NET_84),.T1I2(NET_5),.T1I3(NET_86),.TB1S(GND),.C1Z(NET_204),.Q1Z(m1_ram_control[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_300),.B2I1(m0_m0_control[30]),.B2I2(NET_27),.B2I3(m1_ram_control[30]),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx32122z1),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.B2Z(NET_752),.Q2Z(m1_m1_rnd_dup_0),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M16_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_13_padClk),.QRT(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[5]),.T3I1(lint_ADDR_int[9]),.T3I2(GND),.T3I3(GND),.TB3S(GND),.C3Z(NET_86),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_M17_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000001000),.B0I0(NET_29),.B0I1(NET_34),.B0I2(GND),.B0I3(GND),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_293),.T0I1(m0_coef_wmode_dup_0[1]),.T0I2(m1_m0_dataout_int[11]),.T0I3(NET_66),.TB0S(GND),.B0Z(NET_300),.C0Z(NET_294),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[10]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(i_events[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M17_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_66),.T2I1(m1_ram_control[16]),.T2I2(NET_300),.T2I3(m1_m0_dataout_int[16]),.TB2S(GND),.C2Z(NET_425),.Q2Z(m1_ram_control[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_M17_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx58678z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(m1_m0_dataout_int[10]),.T3I1(NET_63),.T3I2(m0_m1_control[10]),.T3I3(NET_66),.C3Z(NET_272),.Q3Z(m0_m1_control[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_M18_0 (.tFragBitInfo(16'b0000011100000111),.bFragBitInfo(16'b0000000000000111),.B0I0(NET_20),.B0I1(tcdm_result_p0[5]),.B0I2(NET_832),.B0I3(tcdm_result_p2[5]),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(NET_20),.T0I1(tcdm_result_p0[5]),.T0I2(NET_832),.T0I3(tcdm_result_p2[5]),.TB0S(NET_21_CAND4_BLSTR_13_tpGCLKBUF),.C0Z(NET_829),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M18_1 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[5]),.Q1EN(tcdm_valid_p2_int_CAND2_BLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[4]),.T1I1(lint_ADDR_int[3]),.T1I2(lint_ADDR_int[5]),.T1I3(lint_ADDR_int[6]),.TB1S(GND),.C1Z(NET_34),.Q1Z(tcdm_result_p2[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_M18_2 (.tFragBitInfo(16'b0001000100110011),.bFragBitInfo(16'b0000000100000011),.B2I0(NET_300),.B2I1(NET_877),.B2I2(tcdm_result_p2[3]),.B2I3(m1_oper0_wmode_dup_0[1]),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[3]),.Q2EN(tcdm_valid_p2_int_CAND2_BLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T2I0(NET_300),.T2I1(NET_877),.T2I2(tcdm_result_p2[3]),.T2I3(m1_oper0_wmode_dup_0[1]),.TB2S(NET_21_CAND4_BLSTR_13_tpGCLKBUF),.C2Z(NET_874),.Q2Z(tcdm_result_p2[3]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_M18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx10775z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m0_m0_reset_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M19_0 (.tFragBitInfo(16'b0000110011001100),.bFragBitInfo(16'b0000010001000100),.B0I0(tcdm_result_p2[14]),.B0I1(NET_366),.B0I2(tcdm_result_p0[14]),.B0I3(NET_20),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p2[14]),.T0I1(NET_366),.T0I2(tcdm_result_p0[14]),.T0I3(NET_20),.TB0S(NET_21_CAND4_BLSTR_13_tpGCLKBUF),.C0Z(NET_364),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_M19_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[15]),.Q1EN(tcdm_valid_p2_int_CAND2_BLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T1I0(NET_28),.T1I1(fpgaio_in_int[63]),.T1I2(NET_21_CAND4_BLSTR_13_tpGCLKBUF),.T1I3(tcdm_result_p2[31]),.C1Z(NET_776),.Q1Z(tcdm_result_p2[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_M19_2 (.tFragBitInfo(16'b0000011100000111),.bFragBitInfo(16'b0000000000000111),.B2I0(tcdm_result_p0[15]),.B2I1(NET_20),.B2I2(NET_403),.B2I3(tcdm_result_p2[15]),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[14]),.Q2EN(tcdm_valid_p2_int_CAND2_BLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p0[15]),.T2I1(NET_20),.T2I2(NET_403),.T2I3(tcdm_result_p2[15]),.TB2S(NET_21_CAND4_BLSTR_13_tpGCLKBUF),.C2Z(NET_400),.Q2Z(tcdm_result_p2[14]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_M19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_rmode_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[31]),.Q2EN(tcdm_valid_p2_int_CAND2_BLSTR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p2[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M20_3 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'b0000000000000000),.B3I0(NET_8),.B3I1(lint_ADDR_int[14]),.B3I2(lint_ADDR_int[1]),.B3I3(lint_ADDR_int[0]),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[1]),.T3I1(lint_ADDR_int[0]),.T3I2(NET_8),.T3I3(lint_ADDR_int[14]),.TB3S(lint_ADDR_int[10]),.C3Z(NET_5),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_M22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M22_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(GND),.T1I1(lint_ADDR_int[12]),.T1I2(lint_ADDR_int[13]),.T1I3(GND),.TB1S(GND),.C1Z(NET_8),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_M22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[3]),.Q0EN(nx33579z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx33579z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx33579z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx33579z1),.QCK(CLK_int_0__CAND0_BLSTR_13_padClk),.QRT(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_wdata_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[2]),.Q2EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wdata_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_wdata_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdata_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[6]),.Q3EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_waddr_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_M31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[4]),.Q0EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_waddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_M31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[11]),.Q1EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_waddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_M31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[5]),.Q2EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_waddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_M31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[10]),.Q3EN(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_13_padClk),.QRT(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_waddr_dup_0[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[10]),.Q0EN(nx32231z2_CAND4_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_raddr_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[7]),.Q1EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_waddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[0]),.Q2EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_waddr_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[4]),.Q3EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_waddr_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[8]),.Q0EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_waddr_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[9]),.Q1EN(nx32231z2_CAND4_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_raddr_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[11]),.Q2EN(nx32231z2_CAND4_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_raddr_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[8]),.Q3EN(nx32231z2_CAND4_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_raddr_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[5]),.Q0EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_waddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[3]),.Q1EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_waddr_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[9]),.Q2EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_waddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[2]),.Q3EN(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_waddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[0]),.Q3EN(tcdm_valid_p0_int_CAND3_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N5_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_79),.T1I1(NET_78),.T1I2(lint_ADDR_int[12]),.T1I3(GND),.TB1S(GND),.C1Z(nx32231z2),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_N5_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_10),.T2I1(NET_78),.T2I2(lint_ADDR_int[12]),.T2I3(GND),.TB2S(GND),.C2Z(nx15998z1),.Q2Z(m0_coef_we_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[11]),.Q0EN(tcdm_valid_p0_int_CAND3_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[22]),.Q1EN(tcdm_valid_p0_int_CAND3_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[21]),.Q3EN(tcdm_valid_p0_int_CAND3_TLSTR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_14_padClk),.QRT(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[21]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[23]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[23]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N10_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(tcdm_result_p0[0]),.T1I1(NET_126_CAND3_TLSBR_14_tpGCLKBUF),.T1I2(NET_127_CAND4_TLSBR_14_tpGCLKBUF),.T1I3(m0_m1_outsel_dup_0[0]),.C1Z(NET_122),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_N10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000010000),.B0I0(lint_ADDR_int[3]),.B0I1(GND),.B0I2(lint_ADDR_int[2]),.B0I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.B0Z(NET_43),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N11_1 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_25),.T1I1(NET_789),.T1I2(GND),.T1I3(GND),.C1Z(nx50997z2),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_N11_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000001),.B2I0(lint_ADDR_int[3]),.B2I1(GND),.B2I2(lint_ADDR_int[2]),.B2I3(GND),.CD2S(VCC),.Q2DI(lint_WDATA_int[21]),.Q2EN(nx49703z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(tcdm_result_p0[22]),.T2I1(NET_127_CAND4_TLSBR_14_tpGCLKBUF),.T2I2(NET_126_CAND3_TLSBR_14_tpGCLKBUF),.T2I3(m0_m1_control[22]),.TB2S(GND),.B2Z(NET_25),.C2Z(NET_558),.Q2Z(m0_m1_control[21]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_N11_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[22]),.Q3EN(nx49703z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p0[21]),.T3I1(NET_127_CAND4_TLSBR_14_tpGCLKBUF),.T3I2(m0_m1_control[21]),.T3I3(NET_126_CAND3_TLSBR_14_tpGCLKBUF),.C3Z(NET_534),.Q3Z(m0_m1_control[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_N12_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_126_CAND3_TLSBR_14_tpGCLKBUF),.T0I1(NET_127_CAND4_TLSBR_14_tpGCLKBUF),.T0I2(m0_m1_control[23]),.T0I3(tcdm_result_p0[23]),.TB0S(GND),.C0Z(NET_576),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N12_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_24),.T1I1(lint_ADDR_int[11]),.T1I2(NET_4),.T1I3(NET_25),.C1Z(NET_124),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_N12_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_43),.T2I1(lint_ADDR_int[5]),.T2I2(GND),.T2I3(lint_ADDR_int[4]),.TB2S(GND),.C2Z(NET_571),.Q2Z(m0_coef_rmode_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[23]),.Q3EN(nx49703z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_control[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(lint_ADDR_int[3]),.B0I1(lint_ADDR_int[6]),.B0I2(lint_ADDR_int[5]),.B0I3(lint_ADDR_int[4]),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.B0Z(NET_67),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N13_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_207),.T1I1(NET_25),.T1I2(GND),.T1I3(lint_ADDR_int[4]),.TB1S(GND),.Q1Z(m0_m0_clken_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_N13_2 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'b0000000001000000),.B2I0(GND),.B2I1(NET_34),.B2I2(NET_33_CAND2_TLSBR_14_tpGCLKBUF),.B2I3(GND),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(GND),.T2I2(NET_33_CAND2_TLSBR_14_tpGCLKBUF),.T2I3(NET_67),.TB2S(GND),.B2Z(NET_293),.C2Z(NET_65),.Q2Z(m0_ram_control[31]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_N13_3 (.tFragBitInfo(16'b0101111111111111),.bFragBitInfo(16'b0101010101111111),.B3I0(NET_33_CAND2_TLSBR_14_tpGCLKBUF),.B3I1(NET_67),.B3I2(tcdm_wen_p0_dup_0),.B3I3(NET_34),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(tcdm_wen_p0_dup_0),.T3I1(NET_34),.T3I2(NET_33_CAND2_TLSBR_14_tpGCLKBUF),.T3I3(NET_67),.TB3S(m0_ram_control[31]),.C3Z(NET_766),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_N14_0 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b1100100010001000),.B0I0(NET_782),.B0I1(apb_fsm[1]),.B0I2(NET_65),.B0I3(NET_173),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.T0I0(NET_82),.T0I1(lint_ADDR_int[5]),.T0I2(lint_ADDR_int[6]),.T0I3(NET_83),.TB0S(GND),.B0Z(NET_783),.C0Z(NET_207),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N14_1 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.T1I0(NET_33_CAND2_TLSBR_14_tpGCLKBUF),.T1I1(NET_71),.T1I2(GND),.T1I3(GND),.TB1S(GND),.C1Z(NET_241),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_N14_2 (.tFragBitInfo(16'b0111111101111111),.bFragBitInfo(16'b1111111101111111),.B2I0(NET_524),.B2I1(NET_516),.B2I2(NET_921),.B2I3(NET_920),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.T2I0(NET_524),.T2I1(NET_516),.T2I2(NET_921),.T2I3(NET_920),.TB2S(NET_33_CAND2_TLSBR_14_tpGCLKBUF),.Q2Z(lint_RDATA_dup_0[20]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_N14_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.T3I0(NET_82),.T3I1(lint_ADDR_int[9]),.T3I2(NET_4),.T3I3(NET_10),.C3Z(NET_789),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_N15_0 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'b1010101010101000),.B0I0(apb_fsm[0]),.B0I1(NET_78),.B0I2(NET_211),.B0I3(NET_198),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.T0I0(GND),.T0I1(GND),.T0I2(NET_10),.T0I3(lint_ADDR_int[9]),.TB0S(GND),.B0Z(NET_782),.C0Z(NET_83),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N15_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B1I0(NET_925),.B1I1(NET_767),.B1I2(NET_773),.B1I3(NET_771),.CD1S(GND),.Q1DI(GND),.Q1EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.T1I0(NET_773),.T1I1(NET_771),.T1I2(NET_925),.T1I3(NET_767),.TB1S(NET_778),.Q1Z(lint_RDATA_dup_0[31]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_N15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000010000000),.B2I0(NET_5),.B2I1(NET_4),.B2I2(NET_6),.B2I3(lint_ADDR_int[9]),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.B2Z(NET_173),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N15_3 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.T3I0(NET_375),.T3I1(NET_374),.T3I2(NET_377),.T3I3(NET_376),.TB3S(GND),.Q3Z(lint_RDATA_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_N16_0 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0000000000101010),.B0I0(NET_766),.B0I1(NET_300),.B0I2(m1_ram_control[31]),.B0I3(m1_m1_dataout_int[31]),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx49703z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_766),.T0I1(NET_300),.T0I2(m1_ram_control[31]),.T0I3(m1_m1_dataout_int[31]),.TB0S(NET_266),.C0Z(NET_767),.Q0Z(m0_m1_rnd_dup_0),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N16_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(NET_24),.T1I1(NET_22),.T1I2(lint_ADDR_int[11]),.T1I3(NET_4),.C1Z(NET_125),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_N16_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T2I0(NET_84),.T2I1(NET_5),.T2I2(GND),.T2I3(NET_6),.TB2S(GND),.C2Z(NET_82),.Q2Z(m1_ram_control[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_N16_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_0__CAND0_TLSBR_14_padClk),.QRT(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[4]),.T3I1(NET_22),.T3I2(NET_207),.T3I3(GND),.TB3S(GND),.Q3Z(m1_m0_clken_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_N17_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001000000000000),.B0I0(GND),.B0I1(GND),.B0I2(NET_40),.B0I3(NET_33),.T0I0(NET_300),.T0I1(NET_20),.T0I2(tcdm_result_p0[11]),.T0I3(m1_coef_wmode_dup_0[1]),.TB0S(GND),.B0Z(NET_36),.C0Z(NET_298),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_N17_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_299),.T1I1(NET_298),.T1I2(NET_297),.T1I3(NET_296),.C1Z(NET_281),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_N17_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0010000000000000),.B2I0(NET_4),.B2I1(GND),.B2I2(NET_22),.B2I3(NET_24),.T2I0(NET_270),.T2I1(NET_271),.T2I2(NET_272),.T2I3(GND),.TB2S(GND),.B2Z(NET_66),.C2Z(NET_259),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_N17_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_379),.T3I1(NET_378),.T3I2(NET_380),.T3I3(NET_381),.C3Z(NET_375),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_N18_0 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0000010000000000),.B0I0(GND),.B0I1(NET_22),.B0I2(GND),.B0I3(NET_10),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx1800z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T0I0(NET_521),.T0I1(GND),.T0I2(NET_523),.T0I3(NET_522),.TB0S(GND),.B0Z(NET_93),.C0Z(NET_524),.Q0Z(m0_m0_control[20]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_N18_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[9]),.T1I1(NET_82),.T1I2(NET_93),.T1I3(NET_4),.C1Z(nx50995z3),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_N18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000100000000),.B2I0(GND),.B2I1(lint_ADDR_int_2__CAND3_BLSTR_14_tpGCLKBUF),.B2I2(GND),.B2I3(lint_ADDR_int[3]),.CD2S(VCC),.Q2DI(lint_WDATA_int[20]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B2Z(NET_22),.Q2Z(m1_ram_control[20]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N18_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T3I0(NET_27_CAND5_BLSTR_14_tpGCLKBUF),.T3I1(NET_300),.T3I2(m1_ram_control[20]),.T3I3(m0_m0_control[20]),.C3Z(NET_523),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_N19_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_6),.B0I1(NET_5),.B0I2(NET_4),.B0I3(NET_7),.T0I0(lint_ADDR_int[11]),.T0I1(lint_ADDR_int[8]),.T0I2(lint_ADDR_int[9]),.T0I3(GND),.TB0S(GND),.B0Z(NET_2),.C0Z(NET_7),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_N19_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[11]),.T1I1(GND),.T1I2(lint_ADDR_int[7]),.T1I3(lint_ADDR_int[9]),.C1Z(NET_92),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_N19_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_6),.B2I1(NET_5),.B2I2(NET_92),.B2I3(NET_4),.T2I0(NET_93),.T2I1(NET_204),.T2I2(NET_90),.T2I3(GND),.TB2S(GND),.B2Z(NET_90),.C2Z(nx63842z2),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_N19_3 (.tFragBitInfo(16'b0000000100000001),.bFragBitInfo(16'b0000010000000101),.B3I0(NET_2),.B3I1(NET_1),.B3I2(NET_90),.B3I3(NET_204),.T3I0(NET_90),.T3I1(NET_204),.T3I2(NET_2),.T3I3(NET_1),.TB3S(lint_ADDR_int[6]),.C3Z(NET_785),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_N20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N20_2 (.tFragBitInfo(16'b1100110011111111),.bFragBitInfo(16'b0100110001011111),.B2I0(NET_2),.B2I1(tcdm_fmo_p2_int),.B2I2(lint_ADDR_int[7]),.B2I3(tcdm_gnt_p2_int),.T2I0(NET_2),.T2I1(tcdm_fmo_p2_int),.T2I2(lint_ADDR_int[7]),.T2I3(tcdm_gnt_p2_int),.TB2S(NET_93),.C2Z(NET_162),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_N20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_wdsel_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000000000000),.B2I0(lint_ADDR_int[7]),.B2I1(GND),.B2I2(NET_2),.B2I3(NET_93),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B2Z(nx11311z1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N21_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001110111111111),.B3I0(m0_coef_wdsel_dup_0),.B3I1(lint_ADDR_int_2__CAND3_BLSTR_14_tpGCLKBUF),.B3I2(m1_coef_wdsel_dup_0),.B3I3(NET_34),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T3I0(m1_coef_wdsel_dup_0),.T3I1(NET_34),.T3I2(m0_coef_wdsel_dup_0),.T3I3(lint_ADDR_int_2__CAND3_BLSTR_14_tpGCLKBUF),.TB3S(NET_35),.C3Z(NET_366),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_N22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_wdsel_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wmode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000000000000),.B0I0(NET_211),.B0I1(GND),.B0I2(lint_ADDR_int[13]),.B0I3(NET_79),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B0Z(nx14650z1),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N24_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_0__CAND0_BLSTR_14_padClk),.QRT(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF),.QST(GND),.T3I0(NET_211),.T3I1(NET_10),.T3I2(lint_ADDR_int[13]),.T3I3(GND),.TB3S(GND),.C3Z(nx33579z1),.Q3Z(m1_coef_we_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_N26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N26_1 (.tFragBitInfo(16'b0000000000001110),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1EN(nx11311z2),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.T1I0(nx43661z1),.T1I1(nx11311z1),.T1I2(GND),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_req_p2_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.Q1DI(GND),.T1CO());

	LOGIC_2 QL_INST_N26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[1]),.Q0EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_waddr_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[0]),.Q1EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_waddr_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[9]),.Q0EN(nx14650z1_CAND3_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_raddr_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[8]),.Q1EN(nx14650z1_CAND3_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[7]),.Q2EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_waddr_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[2]),.Q3EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_waddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_N31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[3]),.Q0EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_waddr_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_N31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[10]),.Q1EN(nx14650z1_CAND3_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_N31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[9]),.Q2EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_waddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_N31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[8]),.Q3EN(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_14_padClk),.QRT(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_waddr_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[0]),.Q0EN(nx32231z2_CAND4_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q0Z(m0_coef_raddr_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O1_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[1]),.Q1EN(nx32231z2_CAND4_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_raddr_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O1_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[7]),.Q2EN(nx32231z2_CAND4_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_raddr_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[4]),.Q3EN(nx32231z2_CAND4_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_raddr_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O2_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O2_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O2_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[6]),.Q2EN(nx32231z2_CAND4_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_raddr_dup_0[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O2_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[1]),.Q0EN(tcdm_valid_p0_int_CAND3_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[3]),.Q1EN(nx32231z2_CAND4_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q1Z(m0_coef_raddr_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[5]),.Q2EN(nx32231z2_CAND4_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q2Z(m0_coef_raddr_dup_0[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O3_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[2]),.Q3EN(nx32231z2_CAND4_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(m0_coef_raddr_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[9]),.Q3EN(tcdm_valid_p0_int_CAND3_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O6_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m0_m1_dataout_int[16]),.T3I1(fpgaio_in_int[16]),.T3I2(NET_242),.T3I3(NET_69),.TB3S(GND),.C3Z(NET_423),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_O7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[17]),.Q3EN(tcdm_valid_p0_int_CAND3_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[19]),.Q0EN(tcdm_valid_p0_int_CAND3_TLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[19]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_15_padClk),.QRT(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx57183z1),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_outsel_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O10_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(m0_m0_sat_dup_0),.T3I1(NET_107),.T3I2(NET_129),.T3I3(tcdm_addr_p0_dup_0[18]),.TB3S(GND),.C3Z(NET_475),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_O11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[18]),.Q0EN(nx1800z1),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.Q0Z(m0_m0_sat_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O11_1 (.tFragBitInfo(16'b0000110011001100),.bFragBitInfo(16'b0000011100000000),.B1I0(m0_m0_clr_dup_0),.B1I1(NET_129),.B1I2(tcdm_addr_p0_dup_0[17]),.B1I3(NET_442),.CD1S(VCC),.Q1DI(lint_WDATA_int[17]),.Q1EN(nx1800z1),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p0_dup_0[17]),.T1I1(NET_442),.T1I2(m0_m0_clr_dup_0),.T1I3(NET_129),.TB1S(NET_107),.C1Z(NET_439),.Q1Z(m0_m0_clr_dup_0),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_O11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O12_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0010000000000000),.B0I0(NET_24),.B0I1(GND),.B0I2(NET_4),.B0I3(NET_25),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p0[17]),.T0I1(NET_127_CAND4_TLSBR_15_tpGCLKBUF),.T0I2(NET_106),.T0I3(tcdm_result_p2[17]),.TB0S(GND),.B0Z(NET_41),.C0Z(NET_442),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O12_1 (.tFragBitInfo(16'b0111011100000000),.bFragBitInfo(16'b0000010001000100),.B1I0(tcdm_addr_p0_dup_0[19]),.B1I1(NET_490),.B1I2(m0_m0_control[19]),.B1I3(NET_129),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(m0_m0_control[19]),.T1I1(NET_129),.T1I2(tcdm_addr_p0_dup_0[19]),.T1I3(NET_490),.TB1S(NET_107),.C1Z(NET_487),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_O12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000000000000),.B2I0(lint_ADDR_int[11]),.B2I1(NET_23),.B2I2(NET_4),.B2I3(NET_25),.CD2S(VCC),.Q2DI(lint_WDATA_int[19]),.Q2EN(nx1800z1),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.B2Z(NET_127),.Q2Z(m0_m0_control[19]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O12_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p0[19]),.T3I1(NET_127_CAND4_TLSBR_15_tpGCLKBUF),.T3I2(NET_106),.T3I3(tcdm_result_p2[19]),.C3Z(NET_490),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000000000000),.B0I0(GND),.B0I1(NET_23),.B0I2(NET_25),.B0I3(NET_4),.CD0S(VCC),.Q0DI(lint_WDATA_int[16]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.B0Z(NET_20),.Q0Z(m0_ram_control[16]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O13_1 (.tFragBitInfo(16'b0011111100000000),.bFragBitInfo(16'b0000010000001100),.B1I0(m0_m1_dataout_int[31]),.B1I1(NET_924),.B1I2(tcdm_result_p1[31]),.B1I3(NET_69),.CD1S(VCC),.Q1DI(lint_WDATA_int[3]),.Q1EN(nx41096z1),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p1[31]),.T1I1(NET_69),.T1I2(m0_m1_dataout_int[31]),.T1I3(NET_924),.TB1S(NET_42),.C1Z(NET_925),.Q1Z(m1_m1_control[3]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_O13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010001110101111),.B2I0(tcdm_be_p0_dup_0[1]),.B2I1(NET_106),.B2I2(NET_107),.B2I3(tcdm_result_p2[21]),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.B2Z(NET_545),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O13_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p1[16]),.T3I1(m0_ram_control[16]),.T3I2(NET_42),.T3I3(NET_293),.TB3S(GND),.C3Z(NET_420),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_O14_0 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.T0I0(lint_ADDR_int[5]),.T0I1(lint_ADDR_int[4]),.T0I2(lint_ADDR_int[6]),.T0I3(lint_ADDR_int[3]),.TB0S(GND),.C0Z(NET_40),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O14_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.T1I0(NET_424),.T1I1(NET_422),.T1I2(NET_425),.T1I3(NET_423),.C1Z(NET_418),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O14_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_419),.B2I1(NET_420),.B2I2(NET_418),.B2I3(NET_417),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.T2I0(NET_419),.T2I1(NET_420),.T2I2(NET_418),.T2I3(NET_417),.TB2S(NET_421),.Q2Z(lint_RDATA_dup_0[16]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_O14_3 (.tFragBitInfo(16'b1000000010000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_519),.B3I1(tcdm_be_p1_dup_0[0]),.B3I2(NET_520),.B3I3(NET_517),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.T3I0(NET_520),.T3I1(NET_517),.T3I2(NET_519),.T3I3(tcdm_be_p1_dup_0[0]),.TB3S(NET_50),.C3Z(NET_921),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_O15_0 (.tFragBitInfo(16'b0000000000000010),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_42),.B0I1(tcdm_result_p1[4]),.B0I2(NET_37),.B0I3(m1_m1_control[4]),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx41096z1),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T0I0(NET_85),.T0I1(lint_ADDR_int[7]),.T0I2(GND),.T0I3(GND),.TB0S(GND),.B0Z(NET_849),.C0Z(NET_84),.Q0Z(m1_m1_control[4]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O15_1 (.tFragBitInfo(16'b0011000011110000),.bFragBitInfo(16'b0000001000001010),.B1I0(NET_518),.B1I1(tcdm_result_p3[20]),.B1I2(m1_m1_control[20]),.B1I3(NET_64),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_control[20]),.T1I1(NET_64),.T1I2(NET_518),.T1I3(tcdm_result_p3[20]),.TB1S(NET_37),.C1Z(NET_519),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_O15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(m0_m0_dataout_int[31]),.B2I1(NET_64),.B2I2(tcdm_result_p3[31]),.B2I3(NET_41),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.B2Z(NET_768),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0111000000000000),.B3I0(NET_37),.B3I1(m1_m1_reset_dup_0),.B3I2(NET_768),.B3I3(NET_769),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_768),.T3I1(NET_769),.T3I2(NET_37),.T3I3(m1_m1_reset_dup_0),.TB3S(NET_770),.C3Z(NET_771),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_O16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_849),.B0I1(NET_850),.B0I2(NET_851),.B0I3(NET_852),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.B0Z(NET_853),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O16_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.T1I0(NET_331),.T1I1(NET_333),.T1I2(NET_334),.T1I3(NET_332),.C1Z(NET_335),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O16_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_339),.B2I1(NET_342),.B2I2(NET_918),.B2I3(NET_335),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.T2I0(NET_339),.T2I1(NET_342),.T2I2(NET_918),.T2I3(NET_335),.TB2S(NET_349),.Q2Z(lint_RDATA_dup_0[13]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_O16_3 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B3I0(NET_857),.B3I1(NET_928),.B3I2(NET_860),.B3I3(NET_853),.CD3S(GND),.Q3DI(GND),.Q3EN(nx49808z66),.QCK(CLK_int_0__CAND0_TLSBR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF),.T3I0(NET_860),.T3I1(NET_853),.T3I2(NET_857),.T3I3(NET_928),.TB3S(NET_866),.Q3Z(lint_RDATA_dup_0[4]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_O17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_428),.B0I1(NET_427),.B0I2(NET_430),.B0I3(NET_429),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.T0I0(NET_428),.T0I1(NET_427),.T0I2(NET_430),.T0I3(NET_429),.TB0S(NET_431),.C0Z(NET_417),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O17_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.T1I0(NET_27_CAND5_BLSTR_15_tpGCLKBUF),.T1I1(NET_37),.T1I2(m1_m1_rnd_dup_0),.T1I3(m0_m0_rnd_dup_0),.TB1S(GND),.C1Z(NET_430),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_O17_2 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111111111111111),.B2I0(NET_915),.B2I1(NET_245),.B2I2(NET_236),.B2I3(NET_240),.CD2S(GND),.Q2DI(GND),.Q2EN(nx49808z66),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.T2I0(NET_915),.T2I1(NET_245),.T2I2(NET_236),.T2I3(NET_240),.TB2S(NET_252),.Q2Z(lint_RDATA_dup_0[9]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_O17_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.T3I0(NET_234),.T3I1(NET_232),.T3I2(NET_233),.T3I3(NET_235),.TB3S(GND),.C3Z(NET_236),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_O18_0 (.tFragBitInfo(16'b0001000101010101),.bFragBitInfo(16'b0000000100000101),.B0I0(NET_19),.B0I1(NET_20),.B0I2(tcdm_result_p2[1]),.B0I3(tcdm_result_p0[1]),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[19]),.Q0EN(tcdm_valid_p2_int_CAND2_BLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T0I0(NET_19),.T0I1(NET_20),.T0I2(tcdm_result_p2[1]),.T0I3(tcdm_result_p0[1]),.TB0S(NET_21_CAND4_BLSTR_15_tpGCLKBUF),.C0Z(NET_16),.Q0Z(tcdm_result_p2[19]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O18_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[1]),.Q1EN(tcdm_valid_p2_int_CAND2_BLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T1I0(NET_23),.T1I1(lint_ADDR_int[11]),.T1I2(NET_4),.T1I3(NET_22),.C1Z(NET_106),.Q1Z(tcdm_result_p2[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_O18_2 (.tFragBitInfo(16'b0001000101010101),.bFragBitInfo(16'b0000000100000101),.B2I0(NET_237),.B2I1(NET_20),.B2I2(tcdm_result_p2[9]),.B2I3(tcdm_result_p0[9]),.CD2S(VCC),.Q2DI(lint_WDATA_int[16]),.Q2EN(nx1800z1),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_237),.T2I1(NET_20),.T2I2(tcdm_result_p2[9]),.T2I3(tcdm_result_p0[9]),.TB2S(NET_21_CAND4_BLSTR_15_tpGCLKBUF),.C2Z(NET_233),.Q2Z(m0_m0_rnd_dup_0),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_O18_3 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[9]),.Q3EN(tcdm_valid_p2_int_CAND2_BLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_23),.T3I1(GND),.T3I2(NET_4),.T3I3(NET_22),.C3Z(NET_21),.Q3Z(tcdm_result_p2[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[25]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.Q0Z(m0_ram_control[25]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[21]),.Q1EN(tcdm_valid_p2_int_CAND2_BLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O19_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(m0_ram_control[25]),.B2I1(NET_266),.B2I2(NET_293),.B2I3(m1_m1_dataout_int[25]),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T2I0(NET_24),.T2I1(NET_1),.T2I2(m1_m1_dataout_int[9]),.T2I3(NET_4),.TB2S(GND),.B2Z(NET_633),.C2Z(NET_237),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_O19_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T3I0(NET_24),.T3I1(NET_1),.T3I2(m1_m1_dataout_int[1]),.T3I3(NET_4),.C3Z(NET_19),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_O20_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111001101111111),.B0I0(m1_coef_wmode_dup_0[0]),.B0I1(NET_34),.B0I2(lint_ADDR_int_2__CAND3_BLSTR_15_tpGCLKBUF),.B0I3(m0_coef_wmode_dup_0[0]),.CD0S(VCC),.Q0DI(lint_WDATA_int[10]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T0I0(m1_coef_wmode_dup_0[0]),.T0I1(NET_34),.T0I2(lint_ADDR_int_2__CAND3_BLSTR_15_tpGCLKBUF),.T0I3(m0_coef_wmode_dup_0[0]),.TB0S(NET_35),.C0Z(NET_267),.Q0Z(m0_coef_wmode_dup_0[0]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[17]),.Q3EN(tcdm_valid_p2_int_CAND2_BLSTR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p2[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O21_0 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0111001101111111),.B0I0(m1_oper1_rmode_dup_0[1]),.B0I1(NET_34),.B0I2(lint_ADDR_int_2__CAND3_BLSTR_15_tpGCLKBUF),.B0I3(m0_oper1_rmode_dup_0[1]),.CD0S(VCC),.Q0DI(lint_WDATA_int[4]),.Q0EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_rmode_dup_0[1]),.T0I1(NET_34),.T0I2(lint_ADDR_int_2__CAND3_BLSTR_15_tpGCLKBUF),.T0I3(m0_oper1_rmode_dup_0[1]),.TB0S(NET_35),.C0Z(NET_833),.Q0Z(m1_oper1_rmode_dup_0[0]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_O21_1 (.tFragBitInfo(16'b1111111111111111),.bFragBitInfo(16'b0001101111111111),.B1I0(lint_ADDR_int_2__CAND3_BLSTR_15_tpGCLKBUF),.B1I1(m0_oper1_rmode_dup_0[0]),.B1I2(m1_oper1_rmode_dup_0[0]),.B1I3(NET_34),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T1I0(m1_oper1_rmode_dup_0[0]),.T1I1(NET_34),.T1I2(lint_ADDR_int_2__CAND3_BLSTR_15_tpGCLKBUF),.T1I3(m0_oper1_rmode_dup_0[0]),.TB1S(NET_35),.C1Z(NET_855),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_O21_2 (.tFragBitInfo(16'b0101111100000000),.bFragBitInfo(16'b0001001100000000),.B2I0(m0_m0_outsel_dup_0[4]),.B2I1(fpgaio_in_int[36]),.B2I2(NET_27_CAND5_BLSTR_15_tpGCLKBUF),.B2I3(NET_855),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.T2I0(m0_m0_outsel_dup_0[4]),.T2I1(fpgaio_in_int[36]),.T2I2(NET_27_CAND5_BLSTR_15_tpGCLKBUF),.T2I3(NET_855),.TB2S(NET_28),.C2Z(NET_851),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_O21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_wmode_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx49871z1),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.Q2Z(m1_oper1_rmode_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_15_padClk),.QRT(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O26_2 (.tFragBitInfo(16'b0000010100000100),.bFragBitInfo(16'b0000000000000000),.T2I0(GND),.T2I1(p2_fsm[2]),.T2I2(GND),.T2I3(nx11311z1),.TB2S(GND),.C2Z(nx30923z2),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_O26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[0]),.Q0EN(nx14650z1_CAND3_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_raddr_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[1]),.Q2EN(nx14650z1_CAND3_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_raddr_dup_0[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[2]),.Q0EN(nx14650z1_CAND3_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_raddr_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[7]),.Q1EN(nx14650z1_CAND3_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[6]),.Q3EN(nx14650z1_CAND3_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_raddr_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_O31_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_ADDR_int[4]),.Q0EN(nx14650z1_CAND3_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q0Z(m1_coef_raddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_O31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_ADDR_int[11]),.Q1EN(nx14650z1_CAND3_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q1Z(m1_coef_raddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_O31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_ADDR_int[3]),.Q2EN(nx14650z1_CAND3_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q2Z(m1_coef_raddr_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_O31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_ADDR_int[5]),.Q3EN(nx14650z1_CAND3_BLSBR_15_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BLSBR_15_padClk),.QRT(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF),.QST(GND),.Q3Z(m1_coef_raddr_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P4_1 (.tFragBitInfo(16'b0000000000110010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(nx11313z1),.T1I1(GND),.T1I2(p0_fsm[2]),.T1I3(GND),.TB1S(GND),.C1Z(nx41193z2),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_P4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P5_2 (.tFragBitInfo(16'b0000111000000100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.T2I0(nx11313z1),.T2I1(m0_oper0_rdata_int[11]),.T2I2(GND),.T2I3(lint_WDATA_int[11]),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_P5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[16]),.Q3EN(tcdm_valid_p0_int_CAND3_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[31]),.Q3EN(tcdm_valid_p0_int_CAND3_TLSTR_16_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TLSTR_16_padClk),.QRT(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[31]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P9_3 (.tFragBitInfo(16'b0001010101010101),.bFragBitInfo(16'b0000011100001100),.B3I0(m1_coef_rdata_int[11]),.B3I1(lint_ADDR_int[13]),.B3I2(NET_916),.B3I3(lint_ADDR_int[14]),.T3I0(NET_916),.T3I1(lint_ADDR_int[14]),.T3I2(m1_coef_rdata_int[11]),.T3I3(lint_ADDR_int[13]),.TB3S(m0_oper0_rdata_int[11]),.C3Z(NET_929),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_P11_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_3),.B0I1(NET_173),.B0I2(NET_85),.B0I3(NET_43),.T0I0(m0_m0_dataout_int[20]),.T0I1(NET_41),.T0I2(tcdm_result_p1[20]),.T0I3(NET_42),.TB0S(GND),.B0Z(nx11312z1),.C0Z(NET_515),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_P11_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[8]),.T1I1(GND),.T1I2(GND),.T1I3(lint_ADDR_int[11]),.TB1S(GND),.C1Z(NET_85),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_P11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_3),.B2I1(NET_173),.B2I2(NET_85),.B2I3(NET_25),.B2Z(nx11313z1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P11_3 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(GND),.T3I1(NET_789),.T3I2(GND),.T3I3(NET_43),.C3Z(nx50996z2),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[12]),.Q0EN(nx41097z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.Q0Z(m1_m1_mode_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[12]),.Q1EN(nx58678z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_mode_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_P12_2 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(NET_4),.T2I2(NET_43),.T2I3(NET_23),.TB2S(GND),.C2Z(NET_42),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_P12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_P13_0 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(RESET_int[3]),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[5]),.T0I1(lint_ADDR_int[6]),.T0I2(lint_ADDR_int[3]),.T0I3(lint_ADDR_int[4]),.TB0S(GND),.B0Z(not_RESET_3),.C0Z(NET_71),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P13_1 (.tFragBitInfo(16'b0111111101111111),.bFragBitInfo(16'b0001111100111111),.B1I0(m1_m0_control[11]),.B1I1(NET_67),.B1I2(NET_33_CAND2_TLSBR_16_tpGCLKBUF),.B1I3(NET_71),.CD1S(VCC),.Q1DI(lint_WDATA_int[11]),.Q1EN(nx10406z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T1I0(NET_33_CAND2_TLSBR_16_tpGCLKBUF),.T1I1(NET_71),.T1I2(m1_m0_control[11]),.T1I3(NET_67),.TB1S(tcdm_addr_p0_dup_0[11]),.C1Z(NET_291),.Q1Z(m1_m0_control[11]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_P13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_63),.B2I1(NET_41),.B2I2(m0_m1_control[11]),.B2I3(m0_m0_dataout_int[11]),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.B2Z(NET_289),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P13_3 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[11]),.Q3EN(nx58678z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[11]),.T3I1(NET_33_CAND2_TLSBR_16_tpGCLKBUF),.T3I2(GND),.T3I3(NET_67),.C3Z(NET_107),.Q3Z(m0_m1_control[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P14_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000100000),.B0I0(lint_ADDR_int[6]),.B0I1(lint_ADDR_int[4]),.B0I2(lint_ADDR_int[5]),.B0I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(NET_42),.T0I1(NET_37),.T0I2(m1_m1_control[8]),.T0I3(tcdm_result_p1[8]),.TB0S(GND),.B0Z(NET_141),.C0Z(NET_378),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P14_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T1I0(NET_20),.T1I1(NET_64),.T1I2(tcdm_result_p0[16]),.T1I3(tcdm_result_p3[16]),.C1Z(NET_421),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_P14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000010000000),.B2I0(lint_ADDR_int[3]),.B2I1(NET_33_CAND2_TLSBR_16_tpGCLKBUF),.B2I2(NET_141),.B2I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.B2Z(NET_139),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P14_3 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx41097z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_789),.T3I2(GND),.T3I3(NET_1),.C3Z(nx50994z2),.Q3Z(m1_m1_control[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P15_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_4),.T1I1(lint_ADDR_int[11]),.T1I2(NET_1),.T1I3(NET_24),.C1Z(NET_144),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_P15_2 (.tFragBitInfo(16'b0000110011001100),.bFragBitInfo(16'b0000010001000100),.B2I0(tcdm_result_p3[13]),.B2I1(NET_917),.B2I2(m0_m1_dataout_int[13]),.B2I3(NET_69),.T2I0(tcdm_result_p3[13]),.T2I1(NET_917),.T2I2(m0_m1_dataout_int[13]),.T2I3(NET_69),.TB2S(NET_64),.C2Z(NET_918),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_P15_3 (.tFragBitInfo(16'b0011111100000000),.bFragBitInfo(16'b0000010000001100),.B3I0(NET_69),.B3I1(NET_914),.B3I2(tcdm_result_p3[9]),.B3I3(m0_m1_dataout_int[9]),.T3I0(tcdm_result_p3[9]),.T3I1(m0_m1_dataout_int[9]),.T3I2(NET_69),.T3I3(NET_914),.TB3S(NET_64),.C3Z(NET_915),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_P16_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[20]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T0I0(NET_513),.T0I1(NET_515),.T0I2(NET_512),.T0I3(NET_514),.TB0S(GND),.C0Z(NET_516),.Q0Z(m0_ram_control[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P16_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T1I0(NET_4),.T1I1(NET_1),.T1I2(NET_24),.T1I3(GND),.TB1S(GND),.C1Z(NET_266),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_P16_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000001),.B2I0(RESET_int[2]),.B2I1(GND),.B2I2(GND),.B2I3(GND),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T2I0(NET_253),.T2I1(NET_41),.T2I2(tcdm_addr_p2_dup_0[16]),.T2I3(m0_m0_dataout_int[16]),.TB2S(GND),.B2Z(not_RESET_2),.C2Z(NET_424),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_P16_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TLSBR_16_padClk),.QRT(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF),.QST(GND),.T3I0(m0_ram_control[20]),.T3I1(cnt2[1]),.T3I2(NET_36),.T3I3(NET_293),.C3Z(NET_512),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P18_0 (.tFragBitInfo(16'b0000100010001000),.bFragBitInfo(16'b0000000000010000),.B0I0(apb_fsm[0]),.B0I1(GND),.B0I2(lint_ADDR_int[7]),.B0I3(lint_ADDR_int[8]),.T0I0(NET_243),.T0I1(NET_244),.T0I2(fpgaio_oe_dup_0[73]),.T0I3(NET_55),.TB0S(GND),.B0Z(NET_23),.C0Z(NET_245),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_P18_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_776),.T1I1(NET_777),.T1I2(NET_775),.T1I3(NET_774),.C1Z(NET_778),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_P18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(tcdm_result_p0[31]),.B2I1(NET_20),.B2I2(NET_253),.B2I3(tcdm_wen_p2_dup_0),.B2Z(NET_775),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P18_3 (.tFragBitInfo(16'b0100110000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(fpgaio_oe_dup_0[68]),.T3I1(NET_859),.T3I2(NET_55),.T3I3(NET_858),.C3Z(NET_860),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_293),.B0I1(m0_ram_control[27]),.B0I2(m1_m1_dataout_int[27]),.B0I3(NET_266),.CD0S(VCC),.Q0DI(lint_WDATA_int[30]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.B0Z(NET_675),.Q0Z(m0_ram_control[30]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_P19_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T1I0(NET_1),.T1I1(m1_m1_dataout_int[5]),.T1I2(NET_24),.T1I3(NET_4),.C1Z(NET_832),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_P19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001000),.B2I0(lint_ADDR_int_2__CAND3_BLSTR_16_tpGCLKBUF),.B2I1(lint_ADDR_int[3]),.B2I2(GND),.B2I3(GND),.CD2S(VCC),.Q2DI(lint_WDATA_int[27]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.B2Z(NET_1),.Q2Z(m0_ram_control[27]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_P19_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T3I0(NET_293),.T3I1(m0_ram_control[30]),.T3I2(m1_m1_dataout_int[30]),.T3I3(NET_266),.C3Z(NET_747),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_P21_0 (.tFragBitInfo(16'b0000111000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx30923z2),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T0I0(m1_oper0_rdata_int[25]),.T0I1(nx11311z1),.T0I2(GND),.T0I3(lint_WDATA_int[25]),.TB0S(GND),.Q0Z(tcdm_wdata_p2_dup_0[25]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P21_1 (.tFragBitInfo(16'b0000000010111000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx30923z2),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[3]),.T1I1(nx11311z1),.T1I2(m1_oper0_rdata_int[3]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p2_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_P21_2 (.tFragBitInfo(16'b1100111111001111),.bFragBitInfo(16'b1100111110001011),.B2I0(lint_ADDR_int[12]),.B2I1(apb_fsm[0]),.B2I2(lint_ADDR_int[11]),.B2I3(lint_ADDR_int[13]),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[12]),.T2I1(apb_fsm[0]),.T2I2(lint_ADDR_int[11]),.T2I3(lint_ADDR_int[13]),.TB2S(m1_oper0_rdata_int[25]),.C2Z(NET_649),.Q2Z(m0_oper1_rmode_dup_0[0]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_P21_3 (.tFragBitInfo(16'b1100111111001111),.bFragBitInfo(16'b1111110001010101),.B3I0(lint_ADDR_int[11]),.B3I1(lint_ADDR_int[13]),.B3I2(lint_ADDR_int[12]),.B3I3(apb_fsm[0]),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[12]),.T3I1(apb_fsm[0]),.T3I2(lint_ADDR_int[11]),.T3I3(lint_ADDR_int[13]),.TB3S(m1_oper0_rdata_int[3]),.C3Z(NET_886),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_P22_0 (.tFragBitInfo(16'b1111001111110011),.bFragBitInfo(16'b1111001110100011),.B0I0(lint_ADDR_int[12]),.B0I1(lint_ADDR_int[11]),.B0I2(apb_fsm[0]),.B0I3(lint_ADDR_int[13]),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[12]),.T0I1(lint_ADDR_int[11]),.T0I2(apb_fsm[0]),.T0I3(lint_ADDR_int[13]),.TB0S(m1_oper0_rdata_int[10]),.C0Z(NET_276),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_P22_1 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx30923z2),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T1I0(m1_oper0_rdata_int[9]),.T1I1(nx11311z1),.T1I2(lint_WDATA_int[9]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p2_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_P22_2 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx30923z2),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T2I0(nx11311z1),.T2I1(m1_oper0_rdata_int[10]),.T2I2(lint_WDATA_int[10]),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_wdata_p2_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_P22_3 (.tFragBitInfo(16'b1111111100001111),.bFragBitInfo(16'b1101110111010001),.B3I0(lint_ADDR_int[11]),.B3I1(apb_fsm[0]),.B3I2(lint_ADDR_int[12]),.B3I3(lint_ADDR_int[13]),.QCK(CLK_int_0__CAND0_BLSTR_16_padClk),.QRT(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[12]),.T3I1(lint_ADDR_int[13]),.T3I2(lint_ADDR_int[11]),.T3I3(apb_fsm[0]),.TB3S(m1_oper0_rdata_int[9]),.C3Z(NET_247),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_Q4_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.T0I0(m0_coef_rdata_int[22]),.T0I1(m0_oper0_rdata_int[22]),.T0I2(NET_112),.T0I3(NET_61),.TB0S(GND),.C0Z(NET_560),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_Q4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q5_0 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0000000000101010),.B0I0(NET_390),.B0I1(m0_coef_rdata_int[8]),.B0I2(NET_61),.B0I3(m0_oper0_rdata_int[8]),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.T0I0(NET_390),.T0I1(m0_coef_rdata_int[8]),.T0I2(NET_61),.T0I3(m0_oper0_rdata_int[8]),.TB0S(NET_112),.C0Z(NET_389),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[4]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q5_2 (.tFragBitInfo(16'b0101000101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2_CAND3_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(nx11313z1_CAND2_TRSTL_17_tpGCLKBUF),.T2I2(lint_WDATA_int[8]),.T2I3(m0_oper0_rdata_int[8]),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Q5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q6_0 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx41193z2_CAND3_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[22]),.T0I1(GND),.T0I2(nx11313z1_CAND2_TRSTL_17_tpGCLKBUF),.T0I3(m0_oper0_rdata_int[22]),.TB0S(GND),.Q0Z(tcdm_wdata_p0_dup_0[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q6_2 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2_CAND3_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.T2I0(nx11313z1_CAND2_TRSTL_17_tpGCLKBUF),.T2I1(lint_WDATA_int[18]),.T2I2(GND),.T2I3(m0_oper0_rdata_int[18]),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[18]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Q6_3 (.tFragBitInfo(16'b0000111000000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx41193z2_CAND3_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.T3I0(nx11313z1_CAND2_TRSTL_17_tpGCLKBUF),.T3I1(m0_oper0_rdata_int[20]),.T3I2(GND),.T3I3(lint_WDATA_int[20]),.TB3S(GND),.Q3Z(tcdm_wdata_p0_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Q7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[13]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q7_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx41193z2_CAND3_TRSTL_17_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_17_padClk),.QRT(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[25]),.T3I1(m0_oper0_rdata_int[25]),.T3I2(nx11313z1_CAND2_TRSTL_17_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p0_dup_0[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Q9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[25]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[3]),.Q2EN(nx57183z1),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.Q2Z(m0_m1_outsel_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q12_0 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0000000000000000),.T0I0(NET_4),.T0I1(GND),.T0I2(NET_24),.T0I3(NET_43),.TB0S(GND),.C0Z(NET_69),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_Q12_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_oper0_rdata_int[18]),.T1I1(NET_62),.T1I2(m1_oper1_rdata_int[18]),.T1I3(NET_112),.C1Z(NET_464),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Q12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_463),.B2I1(NET_461),.B2I2(NET_462),.B2I3(NET_464),.T2I0(NET_463),.T2I1(NET_461),.T2I2(NET_462),.T2I3(NET_464),.TB2S(NET_465),.C2Z(NET_466),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_Q12_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(tcdm_addr_p0_dup_0[3]),.T3I1(NET_65),.T3I2(NET_37),.T3I3(m1_m1_control[3]),.C3Z(NET_881),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_Q13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_556),.B0I1(NET_557),.B0I2(NET_559),.B0I3(NET_558),.QCK(CLK_int_3__CAND3_TRSBL_17_padClk),.QRT(not_RESET_3),.QST(GND),.T0I0(NET_556),.T0I1(NET_557),.T0I2(NET_559),.T0I3(NET_558),.TB0S(NET_560),.C0Z(NET_552),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q13_1 (.tFragBitInfo(16'b0000000100010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_3__CAND3_TRSBL_17_padClk),.QRT(not_RESET_3),.QST(GND),.T1I0(GND),.T1I1(GND),.T1I2(cnt3[0]),.T1I3(cnt3[1]),.TB1S(GND),.Q1Z(cnt3[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Q13_2 (.tFragBitInfo(16'b0001001000100010),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_457),.B2I1(cnt3[2]),.B2I2(m0_m1_dataout_int[24]),.B2I3(NET_139),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_3__CAND3_TRSBL_17_padClk),.QRT(not_RESET_3),.QST(GND),.T2I0(cnt3[2]),.T2I1(GND),.T2I2(cnt3[0]),.T2I3(cnt3[1]),.TB2S(GND),.B2Z(NET_625),.Q2Z(cnt3[2]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Q13_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_3__CAND3_TRSBL_17_padClk),.QRT(not_RESET_3),.QST(GND),.T3I0(GND),.T3I1(GND),.T3I2(cnt3[0]),.T3I3(GND),.TB3S(GND),.Q3Z(cnt3[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Q14_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B0I0(m1_m0_dataout_int[3]),.B0I1(NET_63),.B0I2(m0_m1_outsel_dup_0[3]),.B0I3(NET_66),.CD0S(VCC),.Q0DI(lint_WDATA_int[8]),.Q0EN(nx10406z1),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T0I0(m1_m0_control[8]),.T0I1(NET_241),.T0I2(m0_m1_control[8]),.T0I3(NET_63),.TB0S(GND),.B0Z(NET_882),.C0Z(NET_392),.Q0Z(m1_m0_control[8]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q14_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T1I0(NET_881),.T1I1(NET_882),.T1I2(GND),.T1I3(NET_880),.C1Z(NET_869),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Q14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Q14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_575),.B3I1(NET_577),.B3I2(NET_576),.B3I3(NET_574),.CD3S(VCC),.Q3DI(lint_WDATA_int[8]),.Q3EN(nx58678z1),.QCK(CLK_int_0__CAND0_TRSBL_17_padClk),.QRT(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF),.QST(GND),.T3I0(NET_576),.T3I1(NET_574),.T3I2(NET_575),.T3I3(NET_577),.TB3S(NET_578),.C3Z(NET_579),.Q3Z(m0_m1_control[8]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Q15_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_36),.B0I1(tcdm_result_p1[30]),.B0I2(cnt5[2]),.B0I3(NET_42),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_5__CAND5_TRSBL_17_padClk),.QRT(not_RESET_2),.QST(GND),.T0I0(GND),.T0I1(cnt5[0]),.T0I2(GND),.T0I3(GND),.TB0S(GND),.B0Z(NET_751),.Q0Z(cnt5[0]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q15_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_5__CAND5_TRSBL_17_padClk),.QRT(not_RESET_2),.QST(GND),.T1I0(NET_139),.T1I1(cnt5[0]),.T1I2(NET_457),.T1I3(m0_m1_dataout_int[28]),.C1Z(NET_706),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Q15_2 (.tFragBitInfo(16'b0001010001010000),.bFragBitInfo(16'b0001001101011111),.B2I0(m0_m1_dataout_int[29]),.B2I1(NET_139),.B2I2(NET_457),.B2I3(cnt5[1]),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_5__CAND5_TRSBL_17_padClk),.QRT(not_RESET_2),.QST(GND),.T2I0(GND),.T2I1(cnt5[0]),.T2I2(cnt5[2]),.T2I3(cnt5[1]),.TB2S(GND),.B2Z(NET_729),.Q2Z(cnt5[2]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Q15_3 (.tFragBitInfo(16'b0000000100000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_5__CAND5_TRSBL_17_padClk),.QRT(not_RESET_2),.QST(GND),.T3I0(GND),.T3I1(cnt5[0]),.T3I2(GND),.T3I3(cnt5[1]),.TB3S(GND),.Q3Z(cnt5[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Q17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100110000000000),.B0I0(NET_55),.B0I1(NET_340),.B0I2(fpgaio_oe_dup_0[77]),.B0I3(NET_341),.B0Z(NET_342),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q17_1 (.tFragBitInfo(16'b0100000011000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_55),.T1I1(NET_884),.T1I2(NET_883),.T1I3(fpgaio_oe_dup_0[67]),.C1Z(NET_880),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Q17_2 (.tFragBitInfo(16'b0111000000000000),.bFragBitInfo(16'b0000011100000000),.B2I0(cnt1[0]),.B2I1(NET_36),.B2I2(GND),.B2I3(NET_426),.T2I0(NET_55),.T2I1(fpgaio_oe_dup_0[74]),.T2I2(NET_273),.T2I3(NET_274),.TB2S(GND),.B2Z(NET_419),.C2Z(NET_270),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_Q17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000010000001100),.B3I0(NET_20),.B3I1(NET_646),.B3I2(NET_645),.B3I3(tcdm_result_p0[25]),.T3I0(NET_645),.T3I1(tcdm_result_p0[25]),.T3I2(NET_20),.T3I3(NET_646),.TB3S(NET_647),.C3Z(NET_644),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_Q18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(tcdm_wen_p3_dup_0),.B0I1(NET_27),.B0I2(NET_70),.B0I3(m0_m0_reset_dup_0),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.B0Z(NET_769),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q18_1 (.tFragBitInfo(16'b0001000100110011),.bFragBitInfo(16'b0000000000010101),.B1I0(tcdm_result_p2[4]),.B1I1(NET_20),.B1I2(tcdm_result_p0[4]),.B1I3(NET_854),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p0[4]),.T1I1(NET_854),.T1I2(tcdm_result_p2[4]),.T1I3(NET_20),.TB1S(NET_21),.C1Z(NET_850),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_Q18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000011000000),.B2I0(fpgaio_oe_dup_0[72]),.B2I1(NET_385),.B2I2(NET_386),.B2I3(NET_55),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_oe_dup_0[72]),.T2I1(NET_385),.T2I2(NET_386),.T2I3(NET_55),.TB2S(NET_387),.C2Z(NET_374),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_Q18_3 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[4]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_728),.T3I2(NET_726),.T3I3(NET_727),.C3Z(NET_723),.Q3Z(tcdm_result_p2[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_Q19_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000001),.B0I0(lint_ADDR_int[8]),.B0I1(GND),.B0I2(apb_fsm_0__CAND4_BRSTL_17_tpGCLKBUF),.B0I3(lint_ADDR_int[7]),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T0I0(m1_m1_dataout_int[16]),.T0I1(NET_28),.T0I2(NET_266),.T0I3(fpgaio_in_int[48]),.TB0S(GND),.B0Z(NET_35),.C0Z(NET_426),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q19_1 (.tFragBitInfo(16'b0000000001110111),.bFragBitInfo(16'b0000000100010001),.B1I0(tcdm_result_p2[13]),.B1I1(NET_336),.B1I2(tcdm_result_p0[13]),.B1I3(NET_20),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[13]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p0[13]),.T1I1(NET_20),.T1I2(tcdm_result_p2[13]),.T1I3(NET_336),.TB1S(NET_21),.C1Z(NET_332),.Q1Z(tcdm_result_p2[13]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_Q19_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T2I0(NET_4),.T2I1(NET_24),.T2I2(m1_m1_dataout_int[15]),.T2I3(NET_1),.TB2S(GND),.C2Z(NET_403),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_Q19_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(RESET_int[0]),.C3Z(not_RESET_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_Q20_0 (.tFragBitInfo(16'b0010001010101010),.bFragBitInfo(16'b0000001000001010),.B0I0(NET_886),.B0I1(m0_coef_rdata_int[3]),.B0I2(m1_oper1_rdata_int[3]),.B0I3(NET_61),.T0I0(NET_886),.T0I1(m0_coef_rdata_int[3]),.T0I2(m1_oper1_rdata_int[3]),.T0I3(NET_61),.TB0S(NET_62_CAND3_BRSTL_17_tpGCLKBUF),.C0Z(NET_883),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_Q20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q20_2 (.tFragBitInfo(16'b0101111100000000),.bFragBitInfo(16'b0001001100000000),.B2I0(m1_oper1_rdata_int[25]),.B2I1(m0_oper0_rdata_int[25]),.B2I2(NET_62_CAND3_BRSTL_17_tpGCLKBUF),.B2I3(NET_649),.T2I0(m1_oper1_rdata_int[25]),.T2I1(m0_oper0_rdata_int[25]),.T2I2(NET_62_CAND3_BRSTL_17_tpGCLKBUF),.T2I3(NET_649),.TB2S(NET_112),.C2Z(NET_646),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_Q20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q21_0 (.tFragBitInfo(16'b0101000011110000),.bFragBitInfo(16'b0001000000110000),.B0I0(NET_62_CAND3_BRSTL_17_tpGCLKBUF),.B0I1(fpgaio_in_int[52]),.B0I2(NET_525),.B0I3(m1_oper1_rdata_int[20]),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T0I0(NET_62_CAND3_BRSTL_17_tpGCLKBUF),.T0I1(fpgaio_in_int[52]),.T0I2(NET_525),.T0I3(m1_oper1_rdata_int[20]),.TB0S(NET_28),.C0Z(NET_522),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q21_1 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T1I0(nx11311z1),.T1I1(lint_WDATA_int[31]),.T1I2(m1_oper0_rdata_int[31]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p2_dup_0[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Q21_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000100010001000),.B2I0(NET_779),.B2I1(NET_780),.B2I2(m1_oper0_rdata_int[31]),.B2I3(NET_113),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T2I0(NET_112),.T2I1(m1_oper0_rdata_int[20]),.T2I2(m0_oper0_rdata_int[20]),.T2I3(NET_113),.TB2S(GND),.B2Z(NET_774),.C2Z(NET_525),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_Q21_3 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T3I0(nx11311z1),.T3I1(GND),.T3I2(lint_WDATA_int[20]),.T3I3(m1_oper0_rdata_int[20]),.TB3S(GND),.Q3Z(tcdm_wdata_p2_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Q22_0 (.tFragBitInfo(16'b0101000001000100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(m1_oper0_rdata_int[8]),.T0I2(lint_WDATA_int[8]),.T0I3(nx11311z1),.TB0S(GND),.Q0Z(tcdm_wdata_p2_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Q22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q22_2 (.tFragBitInfo(16'b0010000010100000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.T2I0(NET_389),.T2I1(m1_oper0_rdata_int[8]),.T2I2(NET_388),.T2I3(NET_113),.TB2S(GND),.C2Z(NET_385),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_Q22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_17_padClk),.QRT(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND2_BRSBL_17_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q25_1 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND2_BRSBL_17_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[22]),.T1I1(m1_oper0_rdata_int[22]),.T1I2(nx11311z1_CAND5_BRSBL_17_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p2_dup_0[22]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Q25_2 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND2_BRSBL_17_tpGCLKBUF),.QST(GND),.T2I0(m1_oper0_rdata_int[23]),.T2I1(lint_WDATA_int[23]),.T2I2(nx11311z1_CAND5_BRSBL_17_tpGCLKBUF),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_wdata_p2_dup_0[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Q25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND2_BRSBL_17_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Q26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND2_BRSBL_17_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q26_1 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND2_BRSBL_17_tpGCLKBUF),.QST(GND),.T1I0(m1_oper0_rdata_int[28]),.T1I1(GND),.T1I2(nx11311z1_CAND5_BRSBL_17_tpGCLKBUF),.T1I3(lint_WDATA_int[28]),.TB1S(GND),.Q1Z(tcdm_wdata_p2_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Q26_2 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND2_BRSBL_17_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[29]),.T2I1(nx11311z1_CAND5_BRSBL_17_tpGCLKBUF),.T2I2(GND),.T2I3(m1_oper0_rdata_int[29]),.TB2S(GND),.Q2Z(tcdm_wdata_p2_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Q26_3 (.tFragBitInfo(16'b0100010001010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_17_padClk),.QRT(not_RESET_0_CAND2_BRSBL_17_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(lint_WDATA_int[18]),.T3I2(m1_oper0_rdata_int[18]),.T3I3(nx11311z1_CAND5_BRSBL_17_tpGCLKBUF),.TB3S(GND),.Q3Z(tcdm_wdata_p2_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Q29_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Q29_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_111),.T2I1(m1_coef_rdata_int[22]),.T2I2(m1_oper0_rdata_int[22]),.T2I3(NET_113_CAND4_BRSBL_17_tpGCLKBUF),.TB2S(GND),.C2Z(NET_559),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_Q29_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_111),.T3I1(NET_113_CAND4_BRSBL_17_tpGCLKBUF),.T3I2(m1_oper0_rdata_int[23]),.T3I3(m1_coef_rdata_int[23]),.C3Z(NET_574),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_Q30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Q30_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m1_oper0_rdata_int[28]),.T1I1(m1_coef_rdata_int[28]),.T1I2(NET_113_CAND4_BRSBL_17_tpGCLKBUF),.T1I3(NET_111),.C1Z(NET_703),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Q30_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_113_CAND4_BRSBL_17_tpGCLKBUF),.B2I1(NET_111),.B2I2(m1_coef_rdata_int[29]),.B2I3(m1_oper0_rdata_int[29]),.T2I0(m1_coef_rdata_int[18]),.T2I1(NET_111),.T2I2(NET_113_CAND4_BRSBL_17_tpGCLKBUF),.T2I3(m1_oper0_rdata_int[18]),.TB2S(GND),.B2Z(NET_726),.C2Z(NET_465),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_Q30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R4_2 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2_CAND3_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T2I0(nx11313z1_CAND2_TRSTL_18_tpGCLKBUF),.T2I1(m0_oper0_rdata_int[4]),.T2I2(lint_WDATA_int[4]),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_R4_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T3I0(m0_coef_rdata_int[21]),.T3I1(m0_oper0_rdata_int[21]),.T3I2(NET_112),.T3I3(NET_61),.C3Z(NET_536),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_R5_0 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx41193z2_CAND3_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[5]),.T0I1(m0_oper0_rdata_int[5]),.T0I2(nx11313z1_CAND2_TRSTL_18_tpGCLKBUF),.T0I3(GND),.TB0S(GND),.Q0Z(tcdm_wdata_p0_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R5_1 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx41193z2_CAND3_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T1I0(nx11313z1_CAND2_TRSTL_18_tpGCLKBUF),.T1I1(m0_oper0_rdata_int[9]),.T1I2(lint_WDATA_int[9]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p0_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_R5_2 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2_CAND3_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T2I0(nx11313z1_CAND2_TRSTL_18_tpGCLKBUF),.T2I1(lint_WDATA_int[15]),.T2I2(GND),.T2I3(m0_oper0_rdata_int[15]),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_R5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p0_int[8]),.Q3EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R6_2 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2_CAND3_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_WDATA_int[21]),.T2I2(nx11313z1_CAND2_TRSTL_18_tpGCLKBUF),.T2I3(m0_oper0_rdata_int[21]),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[21]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_R6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[10]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R7_1 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx41193z2_CAND3_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[31]),.T1I1(m0_oper0_rdata_int[31]),.T1I2(nx11313z1_CAND2_TRSTL_18_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p0_dup_0[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_R7_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[12]),.T2I1(apb_fsm[0]),.T2I2(GND),.T2I3(lint_ADDR_int[13]),.TB2S(GND),.C2Z(NET_61),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_R7_3 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx41193z2_CAND3_TRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_18_padClk),.QRT(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF),.QST(GND),.T3I0(m0_oper0_rdata_int[29]),.T3I1(nx11313z1_CAND2_TRSTL_18_tpGCLKBUF),.T3I2(lint_WDATA_int[29]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p0_dup_0[29]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_R9_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0111101111111011),.B0I0(lint_ADDR_int[13]),.B0I1(apb_fsm[0]),.B0I2(lint_ADDR_int[14]),.B0I3(m1_coef_rdata_int[9]),.T0I0(lint_ADDR_int[13]),.T0I1(apb_fsm[0]),.T0I2(lint_ADDR_int[14]),.T0I3(m1_coef_rdata_int[9]),.TB0S(m0_oper0_rdata_int[9]),.C0Z(NET_246),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_R9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R10_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0111101011111111),.B0I0(lint_ADDR_int[13]),.B0I1(m1_coef_rdata_int[4]),.B0I2(lint_ADDR_int[14]),.B0I3(apb_fsm[0]),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[13]),.T0I1(m1_coef_rdata_int[4]),.T0I2(lint_ADDR_int[14]),.T0I3(apb_fsm[0]),.TB0S(m0_oper0_rdata_int[4]),.C0Z(NET_861),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R10_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0111110011111111),.B2I0(m1_coef_rdata_int[5]),.B2I1(lint_ADDR_int[13]),.B2I2(lint_ADDR_int[14]),.B2I3(apb_fsm[0]),.CD2S(VCC),.Q2DI(lint_WDATA_int[1]),.Q2EN(nx57183z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(m1_coef_rdata_int[5]),.T2I1(lint_ADDR_int[13]),.T2I2(lint_ADDR_int[14]),.T2I3(apb_fsm[0]),.TB2S(m0_oper0_rdata_int[5]),.C2Z(NET_839),.Q2Z(m0_m1_outsel_dup_0[1]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_R10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[5]),.Q3EN(nx57183z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_outsel_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_241),.B0I1(tcdm_addr_p0_dup_0[16]),.B0I2(m1_m0_rnd_dup_0),.B0I3(NET_65),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.B0Z(NET_422),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx10406z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.Q1Z(m1_m0_osel_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[10]),.Q2EN(nx10406z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.Q2Z(m1_m0_control[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R11_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx10406z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T3I0(m0_m1_dataout_int[14]),.T3I1(NET_241),.T3I2(m1_m0_osel_dup_0),.T3I3(NET_69),.TB3S(GND),.C3Z(NET_372),.Q3Z(m1_m0_csel_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_R12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_532),.B0I1(NET_535),.B0I2(NET_533),.B0I3(NET_534),.CD0S(VCC),.Q0DI(lint_WDATA_int[13]),.Q0EN(nx58678z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(NET_532),.T0I1(NET_535),.T0I2(NET_533),.T0I3(NET_534),.TB0S(NET_536),.C0Z(NET_537),.Q0Z(m0_m1_mode_dup_0[1]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000000000000),.B1I0(NET_499),.B1I1(NET_498),.B1I2(NET_496),.B1I3(NET_497),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(NET_496),.T1I1(NET_497),.T1I2(NET_499),.T1I3(NET_498),.TB1S(NET_500),.C1Z(NET_489),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_R12_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[4]),.Q2EN(nx57183z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(NET_241),.T2I1(NET_63),.T2I2(m1_m0_csel_dup_0),.T2I3(m0_m1_csel_dup_0),.TB2S(GND),.C2Z(NET_414),.Q2Z(m0_m1_outsel_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_R12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[15]),.Q3EN(nx58678z1),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.Q3Z(m0_m1_csel_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R13_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(cnt3[0]),.B0I1(NET_145),.B0I2(tcdm_result_p1[22]),.B0I3(NET_139),.T0I0(NET_538),.T0I1(NET_541),.T0I2(NET_540),.T0I3(NET_539),.TB0S(GND),.B0Z(NET_561),.C0Z(NET_542),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_R13_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_562),.T1I1(NET_563),.T1I2(NET_564),.T1I3(NET_561),.C1Z(NET_553),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_R13_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_145),.B2I1(tcdm_result_p1[23]),.B2I2(cnt3[1]),.B2I3(NET_139),.T2I0(tcdm_result_p1[21]),.T2I1(NET_145),.T2I2(cnt2[2]),.T2I3(NET_139),.TB2S(GND),.B2Z(NET_580),.C2Z(NET_538),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_R13_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_581),.T3I1(NET_582),.T3I2(NET_580),.T3I3(NET_583),.C3Z(NET_584),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_R14_0 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_416),.B0I1(NET_414),.B0I2(NET_415),.B0I3(NET_413),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(NET_4),.T0I1(NET_35),.T0I2(NET_43),.T0I3(GND),.TB0S(GND),.B0Z(NET_398),.C0Z(NET_50),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R14_1 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(NET_207),.T1I1(GND),.T1I2(NET_43),.T1I3(lint_ADDR_int[4]),.TB1S(GND),.Q1Z(m0_m1_clken_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_R14_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_241),.B2I1(m1_m0_outsel_dup_0[5]),.B2I2(NET_63),.B2I3(m0_m1_outsel_dup_0[5]),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p0_dup_0[15]),.T2I1(m1_m0_dataout_int[15]),.T2I2(NET_66),.T2I3(NET_65),.TB2S(GND),.B2Z(NET_842),.C2Z(NET_415),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_R14_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_0__CAND0_TRSBL_18_padClk),.QRT(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF),.QST(GND),.T3I0(NET_207),.T3I1(NET_1),.T3I2(lint_ADDR_int[4]),.T3I3(GND),.TB3S(GND),.Q3Z(m1_m1_clken_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_R15_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B0I0(m1_m0_dataout_int[31]),.B0I1(tcdm_wen_p1_dup_0),.B0I2(NET_50),.B0I3(NET_66),.QCK(CLK_int_2__CAND2_TRSBL_18_padClk),.QRT(not_RESET_2),.QST(GND),.T0I0(NET_139),.T0I1(m0_m1_dataout_int[26]),.T0I2(cnt4[1]),.T0I3(NET_457),.TB0S(GND),.B0Z(NET_777),.C0Z(NET_664),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R15_1 (.tFragBitInfo(16'b0001001100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_2__CAND2_TRSBL_18_padClk),.QRT(not_RESET_2),.QST(GND),.T1I0(cnt2[0]),.T1I1(GND),.T1I2(cnt2[1]),.T1I3(cnt2[2]),.TB1S(GND),.Q1Z(cnt2[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_R15_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B2I0(m1_m0_dataout_int[4]),.B2I1(tcdm_addr_p0_dup_0[4]),.B2I2(NET_65),.B2I3(NET_66),.QCK(CLK_int_2__CAND2_TRSBL_18_padClk),.QRT(not_RESET_2),.QST(GND),.T2I0(NET_63),.T2I1(m1_m0_dataout_int[13]),.T2I2(NET_66),.T2I3(m0_m1_mode_dup_0[1]),.TB2S(GND),.B2Z(NET_865),.C2Z(NET_345),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_R15_3 (.tFragBitInfo(16'b0000000100000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_2__CAND2_TRSBL_18_padClk),.QRT(not_RESET_2),.QST(GND),.T3I0(cnt2[0]),.T3I1(GND),.T3I2(GND),.T3I3(cnt2[1]),.TB3S(GND),.Q3Z(cnt2[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_R16_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0001010100111111),.B0I0(tcdm_result_p3[4]),.B0I1(NET_63),.B0I2(m0_m1_outsel_dup_0[4]),.B0I3(NET_64),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_2__CAND2_TRSBL_18_padClk),.QRT(not_RESET_2),.QST(GND),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(cnt2[0]),.TB0S(GND),.B0Z(NET_864),.Q0Z(cnt2[0]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R16_1 (.tFragBitInfo(16'b0000101010101010),.bFragBitInfo(16'b0000000001110000),.B1I0(NET_139),.B1I1(cnt2[0]),.B1I2(NET_501),.B1I3(tcdm_result_p3[19]),.QCK(CLK_int_2__CAND2_TRSBL_18_padClk),.QRT(not_RESET_2),.QST(GND),.T1I0(NET_501),.T1I1(tcdm_result_p3[19]),.T1I2(NET_139),.T1I3(cnt2[0]),.TB1S(NET_140),.C1Z(NET_497),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_R16_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_863),.B2I1(NET_864),.B2I2(GND),.B2I3(NET_865),.QCK(CLK_int_2__CAND2_TRSBL_18_padClk),.QRT(not_RESET_2),.QST(GND),.T2I0(NET_288),.T2I1(NET_286),.T2I2(NET_287),.T2I3(NET_289),.TB2S(GND),.B2Z(NET_866),.C2Z(NET_282),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_R16_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_2__CAND2_TRSBL_18_padClk),.QRT(not_RESET_2),.QST(GND),.T3I0(m0_m1_outsel_dup_0[1]),.T3I1(NET_63),.T3I2(tcdm_result_p3[1]),.T3I3(NET_64),.C3Z(NET_44),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_R17_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[23]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T0I0(m1_m0_dataout_int[14]),.T0I1(NET_63),.T0I2(m0_m1_osel_dup_0),.T0I3(NET_66),.TB0S(GND),.C0Z(NET_362),.Q0Z(m0_ram_control[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx58678z1),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.Q1Z(m0_m1_osel_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R17_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001001101011111),.B2I0(m1_m0_dataout_int[9]),.B2I1(NET_63),.B2I2(NET_66),.B2I3(m0_m1_control[9]),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T2I0(m0_m1_rnd_dup_0),.T2I1(NET_63),.T2I2(tcdm_addr_p3_dup_0[16]),.T2I3(NET_70),.TB2S(GND),.B2Z(NET_248),.C2Z(NET_427),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_R17_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[9]),.Q3EN(nx58678z1),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T3I0(m0_ram_control[23]),.T3I1(NET_140),.T3I2(NET_142),.T3I3(tcdm_result_p3[23]),.TB3S(GND),.C3Z(NET_575),.Q3Z(m0_m1_control[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_R18_0 (.tFragBitInfo(16'b0001000101010101),.bFragBitInfo(16'b0000000100000101),.B0I0(NET_382),.B0I1(NET_20),.B0I2(tcdm_result_p2[8]),.B0I3(tcdm_result_p0[8]),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T0I0(NET_382),.T0I1(NET_20),.T0I2(tcdm_result_p2[8]),.T0I3(tcdm_result_p0[8]),.TB0S(NET_21),.C0Z(NET_379),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R18_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T1I0(NET_266),.T1I1(NET_20),.T1I2(m1_m1_dataout_int[10]),.T1I3(tcdm_result_p0[10]),.C1Z(NET_264),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_R18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R18_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[8]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T3I0(NET_112),.T3I1(NET_62_CAND3_BRSTL_18_tpGCLKBUF),.T3I2(m1_oper1_rdata_int[29]),.T3I3(m0_oper0_rdata_int[29]),.C3Z(NET_728),.Q3Z(tcdm_result_p2[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_R19_0 (.tFragBitInfo(16'b0101111100000000),.bFragBitInfo(16'b0001001100000000),.B0I0(NET_61),.B0I1(m1_oper1_rdata_int[4]),.B0I2(m0_coef_rdata_int[4]),.B0I3(NET_862),.T0I0(NET_61),.T0I1(m1_oper1_rdata_int[4]),.T0I2(m0_coef_rdata_int[4]),.T0I3(NET_862),.TB0S(NET_62_CAND3_BRSTL_18_tpGCLKBUF),.C0Z(NET_858),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_R19_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_24),.T1I1(NET_1),.T1I2(NET_4),.T1I3(m1_m1_dataout_int[3]),.C1Z(NET_877),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_R19_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_703),.B2I1(NET_704),.B2I2(GND),.B2I3(NET_705),.T2I0(m1_m1_dataout_int[13]),.T2I1(NET_24),.T2I2(NET_4),.T2I3(NET_1),.TB2S(GND),.B2Z(NET_700),.C2Z(NET_336),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_R19_3 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(GND),.T3I1(NET_622),.T3I2(NET_623),.T3I3(NET_624),.C3Z(NET_619),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_R20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R20_1 (.tFragBitInfo(16'b0010001010101010),.bFragBitInfo(16'b0001000001010000),.B1I0(m1_oper1_rdata_int[10]),.B1I1(m0_coef_rdata_int[10]),.B1I2(NET_276),.B1I3(NET_61),.T1I0(NET_276),.T1I1(NET_61),.T1I2(m1_oper1_rdata_int[10]),.T1I3(m0_coef_rdata_int[10]),.TB1S(NET_62_CAND3_BRSTL_18_tpGCLKBUF),.C1Z(NET_273),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_R20_2 (.tFragBitInfo(16'b0100010011001100),.bFragBitInfo(16'b0000010000001100),.B2I0(NET_61),.B2I1(NET_344),.B2I2(m1_oper1_rdata_int[13]),.B2I3(m0_coef_rdata_int[13]),.T2I0(NET_61),.T2I1(NET_344),.T2I2(m1_oper1_rdata_int[13]),.T2I3(m0_coef_rdata_int[13]),.TB2S(NET_62_CAND3_BRSTL_18_tpGCLKBUF),.C2Z(NET_340),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_R20_3 (.tFragBitInfo(16'b0101000011110000),.bFragBitInfo(16'b0000000000101010),.B3I0(NET_247),.B3I1(m0_coef_rdata_int[9]),.B3I2(NET_61),.B3I3(m1_oper1_rdata_int[9]),.T3I0(NET_61),.T3I1(m1_oper1_rdata_int[9]),.T3I2(NET_247),.T3I3(m0_coef_rdata_int[9]),.TB3S(NET_62_CAND3_BRSTL_18_tpGCLKBUF),.C3Z(NET_243),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_R21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R21_1 (.tFragBitInfo(16'b1111010111110101),.bFragBitInfo(16'b1010111110001101),.B1I0(apb_fsm_0__CAND4_BRSTL_18_tpGCLKBUF),.B1I1(lint_ADDR_int[12]),.B1I2(lint_ADDR_int[11]),.B1I3(lint_ADDR_int_13__CAND5_BRSTL_18_tpGCLKBUF),.CD1S(VCC),.Q1DI(lint_WDATA_int[5]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[11]),.T1I1(lint_ADDR_int_13__CAND5_BRSTL_18_tpGCLKBUF),.T1I2(apb_fsm_0__CAND4_BRSTL_18_tpGCLKBUF),.T1I3(lint_ADDR_int[12]),.TB1S(m1_oper0_rdata_int[13]),.C1Z(NET_344),.Q1Z(m0_oper1_rmode_dup_0[1]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_R21_2 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[13]),.T2I1(GND),.T2I2(nx11311z1),.T2I3(m1_oper0_rdata_int[13]),.TB2S(GND),.Q2Z(tcdm_wdata_p2_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_R21_3 (.tFragBitInfo(16'b0100010011001100),.bFragBitInfo(16'b0001010100000000),.B3I0(m0_oper0_rdata_int[31]),.B3I1(NET_62_CAND3_BRSTL_18_tpGCLKBUF),.B3I2(m1_oper1_rdata_int[31]),.B3I3(NET_781),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T3I0(m1_oper1_rdata_int[31]),.T3I1(NET_781),.T3I2(m0_oper0_rdata_int[31]),.T3I3(NET_62_CAND3_BRSTL_18_tpGCLKBUF),.TB3S(NET_112),.C3Z(NET_780),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_R22_0 (.tFragBitInfo(16'b1111111100001111),.bFragBitInfo(16'b1110111000001111),.B0I0(lint_ADDR_int[12]),.B0I1(lint_ADDR_int_13__CAND5_BRSTL_18_tpGCLKBUF),.B0I2(lint_ADDR_int[11]),.B0I3(apb_fsm_0__CAND4_BRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[12]),.T0I1(lint_ADDR_int_13__CAND5_BRSTL_18_tpGCLKBUF),.T0I2(lint_ADDR_int[11]),.T0I3(apb_fsm_0__CAND4_BRSTL_18_tpGCLKBUF),.TB0S(m1_oper0_rdata_int[16]),.C0Z(NET_437),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R22_1 (.tFragBitInfo(16'b1111111100001111),.bFragBitInfo(16'b1101110111010001),.B1I0(lint_ADDR_int[11]),.B1I1(apb_fsm_0__CAND4_BRSTL_18_tpGCLKBUF),.B1I2(lint_ADDR_int[12]),.B1I3(lint_ADDR_int_13__CAND5_BRSTL_18_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[12]),.T1I1(lint_ADDR_int_13__CAND5_BRSTL_18_tpGCLKBUF),.T1I2(lint_ADDR_int[11]),.T1I3(apb_fsm_0__CAND4_BRSTL_18_tpGCLKBUF),.TB1S(m1_oper0_rdata_int[4]),.C1Z(NET_862),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_R22_2 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_WDATA_int[16]),.T2I2(nx11311z1),.T2I3(m1_oper0_rdata_int[16]),.TB2S(GND),.Q2Z(tcdm_wdata_p2_dup_0[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_R22_3 (.tFragBitInfo(16'b0101000001000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_18_padClk),.QRT(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(m1_oper0_rdata_int[4]),.T3I2(lint_WDATA_int[4]),.T3I3(nx11311z1),.TB3S(GND),.Q3Z(tcdm_wdata_p2_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_R23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R23_3 (.tFragBitInfo(16'b1111010111110101),.bFragBitInfo(16'b0010011110101111),.B3I0(apb_fsm_0__CAND4_BRSTL_18_tpGCLKBUF),.B3I1(lint_ADDR_int_13__CAND5_BRSTL_18_tpGCLKBUF),.B3I2(lint_ADDR_int[11]),.B3I3(lint_ADDR_int[14]),.T3I0(lint_ADDR_int[11]),.T3I1(lint_ADDR_int[14]),.T3I2(apb_fsm_0__CAND4_BRSTL_18_tpGCLKBUF),.T3I3(lint_ADDR_int_13__CAND5_BRSTL_18_tpGCLKBUF),.TB3S(m1_coef_rdata_int[31]),.C3Z(NET_781),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_R25_0 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND2_BRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(nx11311z1_CAND5_BRSBL_18_tpGCLKBUF),.T0I1(m1_oper0_rdata_int[21]),.T0I2(lint_WDATA_int[21]),.T0I3(GND),.TB0S(GND),.Q0Z(tcdm_wdata_p2_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND2_BRSBL_18_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_R25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND2_BRSBL_18_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND2_BRSBL_18_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R26_0 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND2_BRSBL_18_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(lint_WDATA_int[26]),.T0I2(nx11311z1_CAND5_BRSBL_18_tpGCLKBUF),.T0I3(m1_oper0_rdata_int[26]),.TB0S(GND),.Q0Z(tcdm_wdata_p2_dup_0[26]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_R26_1 (.tFragBitInfo(16'b0101010000000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND2_BRSBL_18_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(m1_oper0_rdata_int[24]),.T1I2(nx11311z1_CAND5_BRSBL_18_tpGCLKBUF),.T1I3(lint_WDATA_int[24]),.TB1S(GND),.Q1Z(tcdm_wdata_p2_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_R26_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND2_BRSBL_18_tpGCLKBUF),.QST(GND),.T2I0(NET_62),.T2I1(m1_oper0_rdata_int[21]),.T2I2(NET_113_CAND4_BRSBL_18_tpGCLKBUF),.T2I3(m1_oper1_rdata_int[21]),.TB2S(GND),.C2Z(NET_535),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_R26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_18_padClk),.QRT(not_RESET_0_CAND2_BRSBL_18_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_R30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_113_CAND4_BRSBL_18_tpGCLKBUF),.B0I1(m1_coef_rdata_int[24]),.B0I2(NET_111),.B0I3(m1_oper0_rdata_int[24]),.B0Z(NET_622),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_R30_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m1_oper0_rdata_int[26]),.T1I1(m1_coef_rdata_int[26]),.T1I2(NET_113_CAND4_BRSBL_18_tpGCLKBUF),.T1I3(NET_111),.TB1S(GND),.C1Z(NET_661),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_R30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_R30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_61),.B0I1(m0_oper1_rdata_int[28]),.B0I2(NET_59_CAND5_TRSTL_19_tpGCLKBUF),.B0I3(m0_coef_rdata_int[28]),.B0Z(NET_704),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S3_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_oper1_rdata_int[31]),.T1I1(NET_61),.T1I2(m0_coef_rdata_int[31]),.T1I3(NET_59_CAND5_TRSTL_19_tpGCLKBUF),.C1Z(NET_779),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S3_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_61),.B2I1(NET_59_CAND5_TRSTL_19_tpGCLKBUF),.B2I2(m0_oper1_rdata_int[29]),.B2I3(m0_coef_rdata_int[29]),.T2I0(m0_coef_rdata_int[26]),.T2I1(m0_oper1_rdata_int[26]),.T2I2(NET_59_CAND5_TRSTL_19_tpGCLKBUF),.T2I3(NET_61),.TB2S(GND),.B2Z(NET_727),.C2Z(NET_662),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S3_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m0_oper1_rdata_int[24]),.T3I1(m0_coef_rdata_int[24]),.T3I2(NET_59_CAND5_TRSTL_19_tpGCLKBUF),.T3I3(NET_61),.C3Z(NET_623),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_S4_0 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx41193z2_CAND3_TRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T0I0(m0_oper0_rdata_int[3]),.T0I1(GND),.T0I2(nx11313z1_CAND2_TRSTL_19_tpGCLKBUF),.T0I3(lint_WDATA_int[3]),.TB0S(GND),.Q0Z(tcdm_wdata_p0_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S4_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx41193z2_CAND3_TRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T1I0(m0_oper0_rdata_int[1]),.T1I1(lint_WDATA_int[1]),.T1I2(nx11313z1_CAND2_TRSTL_19_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p0_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_S4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_S4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S5_0 (.tFragBitInfo(16'b0000111000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx41193z2_CAND3_TRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T0I0(m0_oper0_rdata_int[10]),.T0I1(nx11313z1_CAND2_TRSTL_19_tpGCLKBUF),.T0I2(GND),.T0I3(lint_WDATA_int[10]),.TB0S(GND),.Q0Z(tcdm_wdata_p0_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S5_1 (.tFragBitInfo(16'b0011000011110000),.bFragBitInfo(16'b0000001000001010),.B1I0(NET_412),.B1I1(NET_61),.B1I2(m0_oper0_rdata_int[15]),.B1I3(m0_coef_rdata_int[15]),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T1I0(m0_oper0_rdata_int[15]),.T1I1(m0_coef_rdata_int[15]),.T1I2(NET_412),.T1I3(NET_61),.TB1S(NET_112),.C1Z(NET_409),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_S5_2 (.tFragBitInfo(16'b1111000011111111),.bFragBitInfo(16'b1110000011101111),.B2I0(lint_ADDR_int[14]),.B2I1(lint_ADDR_int[12]),.B2I2(apb_fsm[0]),.B2I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[14]),.T2I1(lint_ADDR_int[12]),.T2I2(apb_fsm[0]),.T2I3(lint_ADDR_int[11]),.TB2S(m0_oper1_rdata_int[15]),.C2Z(NET_412),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_S5_3 (.tFragBitInfo(16'b1111000011111111),.bFragBitInfo(16'b1011101110110001),.B3I0(apb_fsm[0]),.B3I1(lint_ADDR_int[11]),.B3I2(lint_ADDR_int[14]),.B3I3(lint_ADDR_int[12]),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[14]),.T3I1(lint_ADDR_int[12]),.T3I2(apb_fsm[0]),.T3I3(lint_ADDR_int[11]),.TB3S(m0_oper1_rdata_int[8]),.C3Z(NET_390),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_S6_0 (.tFragBitInfo(16'b0101010000010000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx41193z2_CAND3_TRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(nx11313z1_CAND2_TRSTL_19_tpGCLKBUF),.T0I2(m0_oper0_rdata_int[23]),.T0I3(lint_WDATA_int[23]),.TB0S(GND),.Q0Z(tcdm_wdata_p0_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S6_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[20]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S6_2 (.tFragBitInfo(16'b0000111000000010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2_CAND3_TRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(m0_oper0_rdata_int[19]),.T2I1(nx11313z1_CAND2_TRSTL_19_tpGCLKBUF),.T2I2(GND),.T2I3(lint_WDATA_int[19]),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_S6_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T3I0(NET_112),.T3I1(NET_59_CAND5_TRSTL_19_tpGCLKBUF),.T3I2(m0_oper0_rdata_int[23]),.T3I3(m0_oper1_rdata_int[23]),.TB3S(GND),.C3Z(NET_578),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_S7_0 (.tFragBitInfo(16'b0000000000111111),.bFragBitInfo(16'b0000000000010101),.B0I0(m0_oper1_rdata_int[30]),.B0I1(m0_coef_rdata_int[30]),.B0I2(NET_61),.B0I3(NET_762),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T0I0(m0_oper1_rdata_int[30]),.T0I1(m0_coef_rdata_int[30]),.T0I2(NET_61),.T0I3(NET_762),.TB0S(NET_59_CAND5_TRSTL_19_tpGCLKBUF),.C0Z(NET_761),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p0_int[27]),.Q1EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S7_2 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2_CAND3_TRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[27]),.T2I1(m0_oper0_rdata_int[27]),.T2I2(nx11313z1_CAND2_TRSTL_19_tpGCLKBUF),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[27]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_S7_3 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx41193z2_CAND3_TRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.T3I0(m0_oper0_rdata_int[30]),.T3I1(GND),.T3I2(nx11313z1_CAND2_TRSTL_19_tpGCLKBUF),.T3I3(lint_WDATA_int[30]),.TB3S(GND),.Q3Z(tcdm_wdata_p0_dup_0[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_S8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p0_int[30]),.Q0EN(tcdm_valid_p0_int),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_S8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_19_padClk),.QRT(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S9_1 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0111111110111011),.B1I0(lint_ADDR_int[14]),.B1I1(apb_fsm[0]),.B1I2(m1_coef_rdata_int[1]),.B1I3(lint_ADDR_int[13]),.T1I0(m1_coef_rdata_int[1]),.T1I1(lint_ADDR_int[13]),.T1I2(lint_ADDR_int[14]),.T1I3(apb_fsm[0]),.TB1S(m0_oper0_rdata_int[1]),.C1Z(NET_58),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_S9_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0111110111111101),.B2I0(apb_fsm[0]),.B2I1(lint_ADDR_int[13]),.B2I2(lint_ADDR_int[14]),.B2I3(m1_coef_rdata_int[3]),.T2I0(apb_fsm[0]),.T2I1(lint_ADDR_int[13]),.T2I2(lint_ADDR_int[14]),.T2I3(m1_coef_rdata_int[3]),.TB2S(m0_oper0_rdata_int[3]),.C2Z(NET_885),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S9_3 (.tFragBitInfo(16'b0000010000001100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_59),.T3I1(NET_885),.T3I2(GND),.T3I3(m0_oper1_rdata_int[3]),.C3Z(NET_884),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_S10_0 (.tFragBitInfo(16'b0000000000000010),.bFragBitInfo(16'b0000010000001100),.B0I0(m0_oper1_rdata_int[4]),.B0I1(NET_861),.B0I2(GND),.B0I3(NET_59),.T0I0(apb_fsm[0]),.T0I1(lint_ADDR_int[14]),.T0I2(lint_ADDR_int[12]),.T0I3(GND),.TB0S(GND),.B0Z(NET_859),.C0Z(NET_59),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_S10_1 (.tFragBitInfo(16'b0000001000100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_839),.T1I1(GND),.T1I2(m0_oper1_rdata_int[5]),.T1I3(NET_59),.C1Z(NET_838),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S10_2 (.tFragBitInfo(16'b0000000001110111),.bFragBitInfo(16'b0000000000000111),.B2I0(m0_coef_rdata_int[27]),.B2I1(NET_61),.B2I2(m0_oper1_rdata_int[27]),.B2I3(NET_690),.T2I0(m0_coef_rdata_int[27]),.T2I1(NET_61),.T2I2(m0_oper1_rdata_int[27]),.T2I3(NET_690),.TB2S(NET_59),.C2Z(NET_689),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S10_3 (.tFragBitInfo(16'b0000010101010101),.bFragBitInfo(16'b0000000000000111),.B3I0(m0_coef_rdata_int[25]),.B3I1(NET_61),.B3I2(NET_648),.B3I3(m0_oper1_rdata_int[25]),.T3I0(NET_648),.T3I1(m0_oper1_rdata_int[25]),.T3I2(m0_coef_rdata_int[25]),.T3I3(NET_61),.TB3S(NET_59),.C3Z(NET_647),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_S11_0 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0110111111101111),.B0I0(lint_ADDR_int[14]),.B0I1(lint_ADDR_int[13]),.B0I2(apb_fsm[0]),.B0I3(m1_coef_rdata_int[10]),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[14]),.T0I1(lint_ADDR_int[13]),.T0I2(apb_fsm[0]),.T0I3(m1_coef_rdata_int[10]),.TB0S(m0_oper0_rdata_int[10]),.C0Z(NET_275),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S11_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T1I0(m1_m1_csel_dup_0),.T1I1(NET_42),.T1I2(tcdm_result_p1[15]),.T1I3(NET_37),.C1Z(NET_399),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S11_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[15]),.Q2EN(nx41097z1),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T2I0(NET_241),.T2I1(m0_m1_dataout_int[10]),.T2I2(NET_69),.T2I3(m1_m0_control[10]),.TB2S(GND),.C2Z(NET_277),.Q2Z(m1_m1_csel_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_S11_3 (.tFragBitInfo(16'b0000001000100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T3I0(NET_275),.T3I1(GND),.T3I2(NET_59),.T3I3(m0_oper1_rdata_int[10]),.TB3S(GND),.C3Z(NET_274),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_S12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(m0_m1_dataout_int[18]),.B0I1(NET_144),.B0I2(m1_m1_dataout_int[18]),.B0I3(NET_457),.B0Z(NET_462),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S12_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_m1_dataout_int[19]),.T1I1(NET_144),.T1I2(m1_m1_dataout_int[19]),.T1I3(NET_457),.C1Z(NET_498),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S12_2 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_62),.B2I1(m0_oper0_rdata_int[19]),.B2I2(m1_oper1_rdata_int[19]),.B2I3(NET_112),.T2I0(NET_504),.T2I1(NET_502),.T2I2(NET_503),.T2I3(GND),.TB2S(GND),.B2Z(NET_503),.C2Z(NET_500),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S13_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.T0I0(NET_4),.T0I1(NET_43),.T0I2(NET_35),.T0I3(tcdm_addr_p1_dup_0[16]),.TB0S(GND),.C0Z(NET_432),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_S13_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m1_m1_dataout_int[23]),.T1I1(NET_144),.T1I2(m0_m1_dataout_int[23]),.T1I3(NET_457),.TB1S(GND),.C1Z(NET_583),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_S13_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0100000000000000),.B2I0(GND),.B2I1(lint_ADDR_int[14]),.B2I2(lint_ADDR_int[13]),.B2I3(apb_fsm[0]),.T2I0(m0_m1_dataout_int[21]),.T2I1(NET_144),.T2I2(NET_457),.T2I3(m1_m1_dataout_int[21]),.TB2S(GND),.B2Z(NET_111),.C2Z(NET_541),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S13_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m0_m1_dataout_int[22]),.T3I1(NET_144),.T3I2(NET_457),.T3I3(m1_m1_dataout_int[22]),.TB3S(GND),.C3Z(NET_564),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_S14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_841),.B0I1(NET_844),.B0I2(NET_842),.B0I3(NET_843),.B0Z(NET_823),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S14_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m1_m0_outsel_dup_0[3]),.T1I1(NET_241),.T1I2(NET_69),.T1I3(m0_m1_dataout_int[3]),.C1Z(NET_887),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S14_2 (.tFragBitInfo(16'b0010000000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_1),.B2I1(NET_23),.B2I2(lint_ADDR_int[11]),.B2I3(NET_4),.T2I0(apb_fsm[0]),.T2I1(GND),.T2I2(lint_ADDR_int[12]),.T2I3(lint_ADDR_int[14]),.TB2S(GND),.B2Z(NET_140),.C2Z(NET_62),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S14_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(tcdm_addr_p0_dup_0[5]),.T3I1(NET_65),.T3I2(m1_m0_dataout_int[5]),.T3I3(NET_66),.C3Z(NET_843),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_S15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000100000000000),.B0I0(NET_136),.B0I1(NET_135),.B0I2(GND),.B0I3(NET_137),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.B0Z(NET_97),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S15_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[8]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T1I0(NET_66),.T1I1(tcdm_addr_p0_dup_0[1]),.T1I2(m1_m0_dataout_int[1]),.T1I3(NET_65),.TB1S(GND),.C1Z(NET_47),.Q1Z(i_events[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_S15_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_66),.B2I1(m1_m0_dataout_int[8]),.B2I2(NET_65),.B2I3(tcdm_addr_p0_dup_0[8]),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T2I0(NET_393),.T2I1(NET_394),.T2I2(NET_391),.T2I3(NET_392),.TB2S(GND),.B2Z(NET_393),.C2Z(NET_377),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_S15_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_19_padClk),.QRT(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_in_int[8]),.T3I1(NET_51),.T3I2(i_events[8]),.T3I3(NET_242),.TB3S(GND),.C3Z(NET_391),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_S16_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_20),.B0I1(m1_m1_dataout_int[20]),.B0I2(NET_266),.B0I3(tcdm_result_p0[20]),.T0I0(tcdm_result_p2[11]),.T0I1(m0_m1_dataout_int[11]),.T0I2(NET_21),.T0I3(NET_69),.TB0S(GND),.B0Z(NET_513),.C0Z(NET_286),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_S16_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_21),.T1I1(m0_m1_dataout_int[20]),.T1I2(NET_69),.T1I3(tcdm_result_p2[20]),.TB1S(GND),.C1Z(NET_514),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_S16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001100000000),.B2I0(NET_20),.B2I1(NET_687),.B2I2(tcdm_result_p0[27]),.B2I3(NET_688),.T2I0(NET_20),.T2I1(NET_687),.T2I2(tcdm_result_p0[27]),.T2I3(NET_688),.TB2S(NET_689),.C2Z(NET_686),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_46),.B3I1(NET_44),.B3I2(NET_47),.B3I3(NET_45),.T3I0(NET_47),.T3I1(NET_45),.T3I2(NET_46),.T3I3(NET_44),.TB3S(NET_48),.C3Z(NET_13),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_S17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001000001010000),.B0I0(NET_759),.B0I1(NET_20),.B0I2(NET_760),.B0I3(tcdm_result_p0[30]),.T0I0(NET_759),.T0I1(NET_20),.T0I2(NET_760),.T0I3(tcdm_result_p0[30]),.TB0S(NET_761),.C0Z(NET_758),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_S17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000001001100),.B1I0(NET_21),.B1I1(NET_433),.B1I2(tcdm_result_p2[16]),.B1I3(NET_432),.T1I0(tcdm_result_p2[16]),.T1I1(NET_432),.T1I2(NET_21),.T1I3(NET_433),.TB1S(NET_434),.C1Z(NET_431),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_S17_2 (.tFragBitInfo(16'b0000001100110011),.bFragBitInfo(16'b0000000100010001),.B2I0(fpgaio_in_int[75]),.B2I1(NET_290),.B2I2(tcdm_result_p3[11]),.B2I3(NET_64),.T2I0(fpgaio_in_int[75]),.T2I1(NET_290),.T2I2(tcdm_result_p3[11]),.T2I3(NET_64),.TB2S(NET_36),.C2Z(NET_287),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S17_3 (.tFragBitInfo(16'b0010000010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_54),.T3I1(fpgaio_oe_dup_0[65]),.T3I2(NET_56),.T3I3(NET_55),.C3Z(NET_46),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_S18_0 (.tFragBitInfo(16'b0100000011000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_70),.B0I1(NET_242),.B0I2(fpgaio_in_int[5]),.B0I3(tcdm_addr_p3_dup_0[5]),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T0I0(NET_55),.T0I1(NET_410),.T0I2(NET_409),.T0I3(fpgaio_oe_dup_0[79]),.TB0S(GND),.B0Z(NET_841),.C0Z(NET_406),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S18_1 (.tFragBitInfo(16'b0100110000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T1I0(NET_55),.T1I1(NET_838),.T1I2(fpgaio_oe_dup_0[69]),.T1I3(NET_837),.C1Z(NET_836),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S18_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_4),.B2I1(tcdm_result_p3[27]),.B2I2(NET_1),.B2I3(NET_23),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(NET_70),.T2I1(NET_242),.T2I2(fpgaio_in_int[15]),.T2I3(tcdm_addr_p3_dup_0[15]),.TB2S(GND),.B2Z(NET_687),.C2Z(NET_413),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_S18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[11]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p2[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_1),.B0I1(NET_24),.B0I2(m1_m1_dataout_int[4]),.B0I3(NET_4),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.B0Z(NET_854),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S19_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T1I0(NET_112),.T1I1(m1_oper1_rdata_int[28]),.T1I2(m0_oper0_rdata_int[28]),.T1I3(NET_62_CAND3_BRSTL_19_tpGCLKBUF),.C1Z(NET_705),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S19_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0100000000000000),.B2I0(GND),.B2I1(NET_663),.B2I2(NET_661),.B2I3(NET_662),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(NET_1),.T2I1(NET_24),.T2I2(NET_4),.T2I3(m1_m1_dataout_int[8]),.TB2S(GND),.B2Z(NET_658),.C2Z(NET_382),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_S19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[20]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p2[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S20_0 (.tFragBitInfo(16'b1111111100110011),.bFragBitInfo(16'b1111101000110011),.B0I0(lint_ADDR_int[12]),.B0I1(lint_ADDR_int[11]),.B0I2(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.B0I3(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[12]),.T0I1(lint_ADDR_int[11]),.T0I2(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.T0I3(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.TB0S(m1_oper0_rdata_int[30]),.C0Z(NET_763),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S20_1 (.tFragBitInfo(16'b0101010001010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(p2_fsm[4]),.T1I2(nx63842z2),.T1I3(tcdm_req_p2_dup_0),.C1Z(nx60851z2),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S20_2 (.tFragBitInfo(16'b0100110001001100),.bFragBitInfo(16'b0000000001001100),.B2I0(m1_oper1_rdata_int[30]),.B2I1(NET_763),.B2I2(NET_62_CAND3_BRSTL_19_tpGCLKBUF),.B2I3(m0_oper0_rdata_int[30]),.CD2S(VCC),.Q2DI(tcdm_rdata_p2_int[16]),.Q2EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_rdata_int[30]),.T2I1(NET_763),.T2I2(NET_62_CAND3_BRSTL_19_tpGCLKBUF),.T2I3(m0_oper0_rdata_int[30]),.TB2S(NET_112),.C2Z(NET_760),.Q2Z(tcdm_result_p2[16]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_S20_3 (.tFragBitInfo(16'b0011111100000000),.bFragBitInfo(16'b0000010000001100),.B3I0(m0_coef_rdata_int[1]),.B3I1(NET_60),.B3I2(m1_oper1_rdata_int[1]),.B3I3(NET_61),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T3I0(m1_oper1_rdata_int[1]),.T3I1(NET_61),.T3I2(m0_coef_rdata_int[1]),.T3I3(NET_60),.TB3S(NET_62_CAND3_BRSTL_19_tpGCLKBUF),.C3Z(NET_54),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_S21_0 (.tFragBitInfo(16'b1100110011111111),.bFragBitInfo(16'b1100100011111011),.B0I0(lint_ADDR_int[12]),.B0I1(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.B0I2(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.B0I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[12]),.T0I1(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.T0I2(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.T0I3(lint_ADDR_int[11]),.TB0S(m1_oper0_rdata_int[1]),.C0Z(NET_60),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S21_1 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T1I0(nx11311z1),.T1I1(lint_WDATA_int[30]),.T1I2(m1_oper0_rdata_int[30]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p2_dup_0[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_S21_2 (.tFragBitInfo(16'b0011111100000000),.bFragBitInfo(16'b0001010100000000),.B2I0(m0_oper0_rdata_int[27]),.B2I1(m1_oper1_rdata_int[27]),.B2I2(NET_62_CAND3_BRSTL_19_tpGCLKBUF),.B2I3(NET_691),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(m0_oper0_rdata_int[27]),.T2I1(m1_oper1_rdata_int[27]),.T2I2(NET_62_CAND3_BRSTL_19_tpGCLKBUF),.T2I3(NET_691),.TB2S(NET_112),.C2Z(NET_688),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_S21_3 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T3I0(nx11311z1),.T3I1(lint_WDATA_int[1]),.T3I2(m1_oper0_rdata_int[1]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p2_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_S22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000100),.B0I0(lint_ADDR_int[12]),.B0I1(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.B0I2(GND),.B0I3(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.B0Z(NET_113),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S22_2 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(m1_oper0_rdata_int[27]),.T2I1(nx11311z1),.T2I2(lint_WDATA_int[27]),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_wdata_p2_dup_0[27]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_S22_3 (.tFragBitInfo(16'b1100110011111111),.bFragBitInfo(16'b1111101000110011),.B3I0(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.B3I1(lint_ADDR_int[11]),.B3I2(lint_ADDR_int[12]),.B3I3(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[12]),.T3I1(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.T3I2(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.T3I3(lint_ADDR_int[11]),.TB3S(m1_oper0_rdata_int[27]),.C3Z(NET_691),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_S23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S23_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.T1I1(m1_coef_rdata_int[27]),.T1I2(lint_ADDR_int[14]),.T1I3(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.C1Z(NET_690),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_S23_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.B2I1(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.B2I2(m1_coef_rdata_int[30]),.B2I3(lint_ADDR_int[14]),.T2I0(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.T2I1(m1_coef_rdata_int[15]),.T2I2(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.T2I3(lint_ADDR_int[14]),.TB2S(GND),.B2Z(NET_762),.C2Z(NET_411),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_S23_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF),.T3I1(m1_coef_rdata_int[25]),.T3I2(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF),.T3I3(lint_ADDR_int[14]),.C3Z(NET_648),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_S24_0 (.tFragBitInfo(16'b0011001000010000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T0I0(nx11311z1),.T0I1(GND),.T0I2(m1_oper0_rdata_int[15]),.T0I3(lint_WDATA_int[15]),.TB0S(GND),.Q0Z(tcdm_wdata_p2_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_S24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S24_2 (.tFragBitInfo(16'b0001000101010101),.bFragBitInfo(16'b0000000100000101),.B2I0(NET_411),.B2I1(NET_62_CAND3_BRSTL_19_tpGCLKBUF),.B2I2(m1_oper0_rdata_int[15]),.B2I3(m1_oper1_rdata_int[15]),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.T2I0(NET_411),.T2I1(NET_62_CAND3_BRSTL_19_tpGCLKBUF),.T2I2(m1_oper0_rdata_int[15]),.T2I3(m1_oper1_rdata_int[15]),.TB2S(NET_113),.C2Z(NET_410),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_S24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_19_padClk),.QRT(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_19_padClk),.QRT(not_RESET_0_CAND2_BRSBL_19_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S25_1 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_19_padClk),.QRT(not_RESET_0_CAND2_BRSBL_19_tpGCLKBUF),.QST(GND),.T1I0(nx11311z1_CAND5_BRSBL_19_tpGCLKBUF),.T1I1(lint_WDATA_int[11]),.T1I2(m1_oper0_rdata_int[11]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p2_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_S25_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_19_padClk),.QRT(not_RESET_0_CAND2_BRSBL_19_tpGCLKBUF),.QST(GND),.T2I0(NET_62),.T2I1(NET_113_CAND4_BRSBL_19_tpGCLKBUF),.T2I2(m1_oper0_rdata_int[11]),.T2I3(m1_oper1_rdata_int[11]),.TB2S(GND),.C2Z(NET_295),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_S25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_19_padClk),.QRT(not_RESET_0_CAND2_BRSBL_19_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S26_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(m1_oper1_rdata_int[8]),.B0I1(m1_coef_rdata_int[8]),.B0I2(NET_62),.B0I3(NET_111),.QCK(CLK_int_0__CAND0_BRSBL_19_padClk),.QRT(not_RESET_0_CAND2_BRSBL_19_tpGCLKBUF),.QST(GND),.B0Z(NET_388),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S26_1 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_19_padClk),.QRT(not_RESET_0_CAND2_BRSBL_19_tpGCLKBUF),.QST(GND),.T1I0(nx11311z1_CAND5_BRSBL_19_tpGCLKBUF),.T1I1(lint_WDATA_int[19]),.T1I2(m1_oper0_rdata_int[19]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p2_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_S26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_19_padClk),.QRT(not_RESET_0_CAND2_BRSBL_19_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_S26_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_19_padClk),.QRT(not_RESET_0_CAND2_BRSBL_19_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_S30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_S30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_S30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_S30_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_113_CAND4_BRSBL_19_tpGCLKBUF),.T3I1(NET_111),.T3I2(m1_oper0_rdata_int[19]),.T3I3(m1_coef_rdata_int[19]),.TB3S(GND),.C3Z(NET_502),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_T3_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.T0I0(NET_61),.T0I1(m0_oper1_rdata_int[19]),.T0I2(NET_59_CAND5_TRSTL_20_tpGCLKBUF),.T0I3(m0_coef_rdata_int[19]),.TB0S(GND),.C0Z(NET_504),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_T3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T3_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.T2I0(m0_oper1_rdata_int[18]),.T2I1(NET_61),.T2I2(NET_59_CAND5_TRSTL_20_tpGCLKBUF),.T2I3(m0_coef_rdata_int[18]),.TB2S(GND),.C2Z(NET_461),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_T3_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m0_coef_rdata_int[17]),.T3I1(m0_oper1_rdata_int[17]),.T3I2(NET_59_CAND5_TRSTL_20_tpGCLKBUF),.T3I3(NET_61),.TB3S(GND),.C3Z(NET_456),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_T4_0 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx41193z2_CAND3_TRSTL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T0I0(m0_oper0_rdata_int[0]),.T0I1(nx11313z1_CAND2_TRSTL_20_tpGCLKBUF),.T0I2(lint_WDATA_int[0]),.T0I3(GND),.TB0S(GND),.Q0Z(tcdm_wdata_p0_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T4_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T1I0(m0_oper0_rdata_int[0]),.T1I1(m0_oper1_rdata_int[0]),.T1I2(NET_59_CAND5_TRSTL_20_tpGCLKBUF),.T1I3(NET_112),.C1Z(NET_110),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_T4_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T2I0(m0_oper1_rdata_int[7]),.T2I1(m0_oper0_rdata_int[7]),.T2I2(NET_59_CAND5_TRSTL_20_tpGCLKBUF),.T2I3(NET_112),.TB2S(GND),.C2Z(NET_602),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_T4_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx41193z2_CAND3_TRSTL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[7]),.T3I1(m0_oper0_rdata_int[7]),.T3I2(nx11313z1_CAND2_TRSTL_20_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p0_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_T6_0 (.tFragBitInfo(16'b0000111000000100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx41193z2_CAND3_TRSTL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T0I0(nx11313z1_CAND2_TRSTL_20_tpGCLKBUF),.T0I1(m0_oper0_rdata_int[16]),.T0I2(GND),.T0I3(lint_WDATA_int[16]),.TB0S(GND),.Q0Z(tcdm_wdata_p0_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T6_1 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx41193z2_CAND3_TRSTL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(lint_WDATA_int[13]),.T1I2(nx11313z1_CAND2_TRSTL_20_tpGCLKBUF),.T1I3(m0_oper0_rdata_int[13]),.TB1S(GND),.Q1Z(tcdm_wdata_p0_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_T6_2 (.tFragBitInfo(16'b0010101000101010),.bFragBitInfo(16'b0000000000101010),.B2I0(NET_437),.B2I1(m0_oper0_rdata_int[16]),.B2I2(NET_112),.B2I3(m0_oper1_rdata_int[16]),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T2I0(NET_437),.T2I1(m0_oper0_rdata_int[16]),.T2I2(NET_112),.T2I3(m0_oper1_rdata_int[16]),.TB2S(NET_59_CAND5_TRSTL_20_tpGCLKBUF),.C2Z(NET_433),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_T6_3 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx41193z2_CAND3_TRSTL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T3I0(nx11313z1_CAND2_TRSTL_20_tpGCLKBUF),.T3I1(lint_WDATA_int[14]),.T3I2(m0_oper0_rdata_int[14]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p0_dup_0[14]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_T7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(m0_coef_rdata_int[16]),.B0I1(lint_ADDR_int[12]),.B0I2(lint_ADDR_int[13]),.B0I3(apb_fsm[0]),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.B0Z(NET_435),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T7_1 (.tFragBitInfo(16'b1111000011111111),.bFragBitInfo(16'b0001101110111011),.B1I0(apb_fsm[0]),.B1I1(lint_ADDR_int[11]),.B1I2(lint_ADDR_int[13]),.B1I3(lint_ADDR_int[12]),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[13]),.T1I1(lint_ADDR_int[12]),.T1I2(apb_fsm[0]),.T1I3(lint_ADDR_int[11]),.TB1S(m0_coef_rdata_int[20]),.C1Z(NET_528),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_T7_2 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2_CAND3_TRSTL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_WDATA_int[28]),.T2I2(nx11313z1_CAND2_TRSTL_20_tpGCLKBUF),.T2I3(m0_oper0_rdata_int[28]),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_T7_3 (.tFragBitInfo(16'b0000000000001100),.bFragBitInfo(16'b1011000110100000),.B3I0(lint_ADDR_int[12]),.B3I1(lint_ADDR_int[14]),.B3I2(lint_ADDR_int[13]),.B3I3(m0_oper1_rdata_int[11]),.QCK(CLK_int_0__CAND0_TRSTL_20_padClk),.QRT(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[13]),.T3I1(m0_oper1_rdata_int[11]),.T3I2(lint_ADDR_int[12]),.T3I3(lint_ADDR_int[14]),.TB3S(m0_coef_rdata_int[11]),.C3Z(NET_916),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_T8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000100),.B0I0(lint_ADDR_int[14]),.B0I1(apb_fsm[0]),.B0I2(GND),.B0I3(lint_ADDR_int[13]),.B0Z(NET_112),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_T8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_T9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T9_1 (.tFragBitInfo(16'b0000000001110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_oper1_rdata_int[9]),.T1I1(NET_59),.T1I2(NET_246),.T1I3(GND),.TB1S(GND),.C1Z(NET_244),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_T9_2 (.tFragBitInfo(16'b0000001000001010),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_58),.T2I1(NET_59),.T2I2(GND),.T2I3(m0_oper1_rdata_int[1]),.TB2S(GND),.C2Z(NET_56),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_T9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_T10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T10_2 (.tFragBitInfo(16'b0111111111111111),.bFragBitInfo(16'b0110111111101111),.B2I0(lint_ADDR_int[14]),.B2I1(lint_ADDR_int[13]),.B2I2(apb_fsm[0]),.B2I3(m1_coef_rdata_int[13]),.T2I0(lint_ADDR_int[14]),.T2I1(lint_ADDR_int[13]),.T2I2(apb_fsm[0]),.T2I3(m1_coef_rdata_int[13]),.TB2S(m0_oper0_rdata_int[13]),.C2Z(NET_343),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_T10_3 (.tFragBitInfo(16'b0000000000101010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_343),.T3I1(NET_59),.T3I2(m0_oper1_rdata_int[13]),.T3I3(GND),.TB3S(GND),.C3Z(NET_341),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_T11_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0010101000000000),.B0I0(NET_367),.B0I1(m0_oper1_rdata_int[14]),.B0I2(NET_59),.B0I3(NET_368),.T0I0(m1_coef_rdata_int[14]),.T0I1(NET_112),.T0I2(m0_oper0_rdata_int[14]),.T0I3(NET_111),.TB0S(GND),.B0Z(NET_365),.C0Z(NET_367),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_T11_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_600),.T1I1(NET_602),.T1I2(NET_601),.T1I3(GND),.TB1S(GND),.C1Z(NET_595),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_T11_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B2I0(m1_coef_rdata_int[7]),.B2I1(NET_61),.B2I2(m0_coef_rdata_int[7]),.B2I3(NET_111),.T2I0(NET_111),.T2I1(m1_coef_rdata_int[21]),.T2I2(NET_59),.T2I3(m0_oper1_rdata_int[21]),.TB2S(GND),.B2Z(NET_601),.C2Z(NET_532),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_T11_3 (.tFragBitInfo(16'b0100010011001100),.bFragBitInfo(16'b0001010100000000),.B3I0(m0_oper1_rdata_int[20]),.B3I1(NET_111),.B3I2(m1_coef_rdata_int[20]),.B3I3(NET_528),.T3I0(m1_coef_rdata_int[20]),.T3I1(NET_528),.T3I2(m0_oper1_rdata_int[20]),.T3I3(NET_111),.TB3S(NET_59),.C3Z(NET_527),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_T12_0 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_116),.B0I1(NET_24),.B0I2(m0_m1_dataout_int[12]),.B0I3(NET_4),.T0I0(GND),.T0I1(NET_454),.T0I2(NET_456),.T0I3(NET_455),.TB0S(GND),.B0Z(NET_325),.C0Z(NET_452),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_T12_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m1_m1_dataout_int[17]),.T1I1(NET_457),.T1I2(m0_m1_dataout_int[17]),.T1I3(NET_144),.C1Z(NET_450),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_T12_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000100000000000),.B2I0(NET_116),.B2I1(NET_23),.B2I2(GND),.B2I3(NET_4),.T2I0(NET_116),.T2I1(NET_24),.T2I2(GND),.T2I3(NET_4),.TB2S(GND),.B2Z(NET_145),.C2Z(NET_457),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_T12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000000000000),.B3I0(NET_450),.B3I1(NET_451),.B3I2(NET_448),.B3I3(NET_449),.T3I0(NET_448),.T3I1(NET_449),.T3I2(NET_450),.T3I3(NET_451),.TB3S(NET_452),.C3Z(NET_441),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_T14_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_61),.B0I1(m0_coef_rdata_int[6]),.B0I2(NET_111),.B0I3(m1_coef_rdata_int[6]),.T0I0(NET_61),.T0I1(m0_coef_rdata_int[23]),.T0I2(m1_oper1_rdata_int[23]),.T0I3(NET_62),.TB0S(GND),.B0Z(NET_802),.C0Z(NET_577),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_T14_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_888),.T1I1(NET_887),.T1I2(NET_889),.T1I3(NET_890),.C1Z(NET_872),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_T14_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B2I0(m0_m1_dataout_int[5]),.B2I1(NET_69),.B2I2(NET_64),.B2I3(tcdm_result_p3[5]),.T2I0(tcdm_result_p3[15]),.T2I1(NET_69),.T2I2(NET_64),.T2I3(m0_m1_dataout_int[15]),.TB2S(GND),.B2Z(NET_844),.C2Z(NET_416),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_T14_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_242),.T3I1(fpgaio_in_int[3]),.T3I2(NET_64),.T3I3(tcdm_result_p3[3]),.C3Z(NET_890),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_T15_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_61),.B0I1(m0_coef_rdata_int[2]),.B0I2(m1_coef_rdata_int[2]),.B0I3(NET_111),.T0I0(NET_61),.T0I1(m0_coef_rdata_int[12]),.T0I2(m1_coef_rdata_int[12]),.T0I3(NET_111),.TB0S(GND),.B0Z(NET_903),.C0Z(NET_316),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_T15_1 (.tFragBitInfo(16'b0000001100001111),.bFragBitInfo(16'b0000000100000101),.B1I0(NET_325),.B1I1(NET_139),.B1I2(tcdm_result_p3[12]),.B1I3(fpgaio_in_int[76]),.T1I0(tcdm_result_p3[12]),.T1I1(fpgaio_in_int[76]),.T1I2(NET_325),.T1I3(NET_139),.TB1S(NET_140),.C1Z(NET_323),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_T15_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0100000000000000),.B2I0(GND),.B2I1(NET_110),.B2I2(NET_108),.B2I3(NET_109),.T2I0(NET_69),.T2I1(tcdm_result_p3[8]),.T2I2(NET_64),.T2I3(m0_m1_dataout_int[8]),.TB2S(GND),.B2Z(NET_99),.C2Z(NET_394),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_T15_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_61),.T3I1(m0_coef_rdata_int[0]),.T3I2(m1_coef_rdata_int[0]),.T3I3(NET_111),.C3Z(NET_109),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_T16_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000011101110111),.B0I0(cnt4[0]),.B0I1(NET_36),.B0I2(NET_42),.B0I3(tcdm_result_p1[25]),.CD0S(GND),.Q0DI(GND),.Q0EN(VCC),.QCK(CLK_int_4__CAND4_TRSBL_20_padClk),.QRT(not_RESET_1),.QST(GND),.T0I0(GND),.T0I1(cnt4[0]),.T0I2(GND),.T0I3(GND),.TB0S(GND),.B0Z(NET_637),.Q0Z(cnt4[0]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T16_1 (.tFragBitInfo(16'b0000000000010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(VCC),.QCK(CLK_int_4__CAND4_TRSBL_20_padClk),.QRT(not_RESET_1),.QST(GND),.T1I0(GND),.T1I1(cnt4[0]),.T1I2(cnt4[1]),.T1I3(GND),.TB1S(GND),.Q1Z(cnt4[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_T16_2 (.tFragBitInfo(16'b0000000001101010),.bFragBitInfo(16'b0000011101110111),.B2I0(cnt4[2]),.B2I1(NET_36),.B2I2(NET_42),.B2I3(tcdm_result_p1[27]),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_4__CAND4_TRSBL_20_padClk),.QRT(not_RESET_1),.QST(GND),.T2I0(cnt4[2]),.T2I1(cnt4[0]),.T2I2(cnt4[1]),.T2I3(GND),.TB2S(GND),.B2Z(NET_679),.Q2Z(cnt4[2]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_T16_3 (.tFragBitInfo(16'b0011000011110000),.bFragBitInfo(16'b0000001000001010),.B3I0(NET_291),.B3I1(fpgaio_out_dup_0[75]),.B3I2(tcdm_result_p1[11]),.B3I3(NET_254),.QCK(CLK_int_4__CAND4_TRSBL_20_padClk),.QRT(not_RESET_1),.QST(GND),.T3I0(tcdm_result_p1[11]),.T3I1(NET_254),.T3I2(NET_291),.T3I3(fpgaio_out_dup_0[75]),.TB3S(NET_42),.C3Z(NET_288),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_T17_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0100000000000000),.B0I0(GND),.B0I1(NET_1),.B0I2(NET_4),.B0I3(NET_23),.QCK(CLK_int_1__CAND1_BRSTL_20_padClk),.QRT(not_RESET_1),.QST(GND),.T0I0(NET_277),.T0I1(NET_279),.T0I2(NET_278),.T0I3(NET_280),.TB0S(GND),.B0Z(NET_64),.C0Z(NET_262),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_361),.B1I1(NET_359),.B1I2(NET_360),.B1I3(NET_358),.QCK(CLK_int_1__CAND1_BRSTL_20_padClk),.QRT(not_RESET_1),.QST(GND),.T1I0(NET_360),.T1I1(NET_358),.T1I2(NET_361),.T1I3(NET_359),.TB1S(NET_362),.C1Z(NET_354),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_T17_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0001001101011111),.B2I0(tcdm_result_p3[14]),.B2I1(fpgaio_in_int[14]),.B2I2(NET_64),.B2I3(NET_242),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_1__CAND1_BRSTL_20_padClk),.QRT(not_RESET_1),.QST(GND),.T2I0(cnt1[0]),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(NET_361),.Q2Z(cnt1[0]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_T17_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_1__CAND1_BRSTL_20_padClk),.QRT(not_RESET_1),.QST(GND),.T3I0(tcdm_result_p3[10]),.T3I1(NET_64),.T3I2(fpgaio_in_int[10]),.T3I3(NET_242),.C3Z(NET_280),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_T18_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.T0I0(NET_70),.T0I1(tcdm_addr_p3_dup_0[8]),.T0I2(NET_254),.T0I3(fpgaio_out_dup_0[72]),.TB0S(GND),.C0Z(NET_387),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T18_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p3[30]),.T1I1(NET_1),.T1I2(NET_23),.T1I3(NET_4),.C1Z(NET_759),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_T18_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_23),.B2I1(NET_1),.B2I2(tcdm_result_p3[25]),.B2I3(NET_4),.CD2S(VCC),.Q2DI(lint_WDATA_int[14]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.T2I0(NET_70),.T2I1(tcdm_addr_p3_dup_0[10]),.T2I2(NET_254),.T2I3(fpgaio_out_dup_0[74]),.TB2S(GND),.B2Z(NET_645),.C2Z(NET_279),.Q2Z(i_events[14]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_T18_3 (.tFragBitInfo(16'b0000000001110111),.bFragBitInfo(16'b0000000100010001),.B3I0(i_events[14]),.B3I1(NET_363),.B3I2(fpgaio_out_dup_0[78]),.B3I3(NET_254),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.T3I0(fpgaio_out_dup_0[78]),.T3I1(NET_254),.T3I2(i_events[14]),.T3I3(NET_363),.TB3S(NET_51),.C3Z(NET_359),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_T19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_T19_3 (.tFragBitInfo(16'b0000000000000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int[7]),.T3I1(lint_ADDR_int[8]),.T3I2(apb_fsm_0__CAND4_BRSTL_20_tpGCLKBUF),.T3I3(GND),.C3Z(NET_24),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_T20_0 (.tFragBitInfo(16'b0101111100000000),.bFragBitInfo(16'b0001001100000000),.B0I0(m0_coef_rdata_int[5]),.B0I1(m1_oper1_rdata_int[5]),.B0I2(NET_61),.B0I3(NET_840),.T0I0(m0_coef_rdata_int[5]),.T0I1(m1_oper1_rdata_int[5]),.T0I2(NET_61),.T0I3(NET_840),.TB0S(NET_62_CAND3_BRSTL_20_tpGCLKBUF),.C0Z(NET_837),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_T20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T20_2 (.tFragBitInfo(16'b0000101010101010),.bFragBitInfo(16'b0000001000100010),.B2I0(NET_369),.B2I1(m1_oper1_rdata_int[14]),.B2I2(NET_61),.B2I3(m0_coef_rdata_int[14]),.T2I0(NET_369),.T2I1(m1_oper1_rdata_int[14]),.T2I2(NET_61),.T2I3(m0_coef_rdata_int[14]),.TB2S(NET_62_CAND3_BRSTL_20_tpGCLKBUF),.C2Z(NET_368),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_T20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_T22_0 (.tFragBitInfo(16'b0000110000001010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.T0I0(m1_oper0_rdata_int[14]),.T0I1(lint_WDATA_int[14]),.T0I2(GND),.T0I3(nx11311z1),.TB0S(GND),.Q0Z(tcdm_wdata_p2_dup_0[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T22_1 (.tFragBitInfo(16'b1111001111110011),.bFragBitInfo(16'b1010100011111101),.B1I0(apb_fsm_0__CAND4_BRSTL_20_tpGCLKBUF),.B1I1(lint_ADDR_int_13__CAND5_BRSTL_20_tpGCLKBUF),.B1I2(lint_ADDR_int[12]),.B1I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[12]),.T1I1(lint_ADDR_int[11]),.T1I2(apb_fsm_0__CAND4_BRSTL_20_tpGCLKBUF),.T1I3(lint_ADDR_int_13__CAND5_BRSTL_20_tpGCLKBUF),.TB1S(m1_oper0_rdata_int[5]),.C1Z(NET_840),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_T22_2 (.tFragBitInfo(16'b1111001111110011),.bFragBitInfo(16'b1111001110100011),.B2I0(lint_ADDR_int[12]),.B2I1(lint_ADDR_int[11]),.B2I2(apb_fsm_0__CAND4_BRSTL_20_tpGCLKBUF),.B2I3(lint_ADDR_int_13__CAND5_BRSTL_20_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[12]),.T2I1(lint_ADDR_int[11]),.T2I2(apb_fsm_0__CAND4_BRSTL_20_tpGCLKBUF),.T2I3(lint_ADDR_int_13__CAND5_BRSTL_20_tpGCLKBUF),.TB2S(m1_oper0_rdata_int[14]),.C2Z(NET_369),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_T22_3 (.tFragBitInfo(16'b0000101000001100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[5]),.T3I1(m1_oper0_rdata_int[5]),.T3I2(GND),.T3I3(nx11311z1),.TB3S(GND),.Q3Z(tcdm_wdata_p2_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_T23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T23_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[14]),.T1I1(apb_fsm_0__CAND4_BRSTL_20_tpGCLKBUF),.T1I2(lint_ADDR_int_13__CAND5_BRSTL_20_tpGCLKBUF),.T1I3(m1_coef_rdata_int[16]),.TB1S(GND),.C1Z(NET_436),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_T23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000010101),.B2I0(NET_435),.B2I1(m1_oper1_rdata_int[16]),.B2I2(NET_62_CAND3_BRSTL_20_tpGCLKBUF),.B2I3(NET_436),.B2Z(NET_434),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_T23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_T24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T24_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.T1I0(NET_62_CAND3_BRSTL_20_tpGCLKBUF),.T1I1(NET_113),.T1I2(m1_oper0_rdata_int[7]),.T1I3(m1_oper1_rdata_int[7]),.TB1S(GND),.C1Z(NET_600),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_T24_2 (.tFragBitInfo(16'b0000000010111000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[7]),.T2I1(nx11311z1),.T2I2(m1_oper0_rdata_int[7]),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_wdata_p2_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_T24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_20_padClk),.QRT(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_T25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_62),.B0I1(m1_oper1_rdata_int[2]),.B0I2(NET_113_CAND4_BRSBL_20_tpGCLKBUF),.B0I3(m1_oper0_rdata_int[2]),.QCK(CLK_int_0__CAND0_BRSBL_20_padClk),.QRT(not_RESET_0_CAND2_BRSBL_20_tpGCLKBUF),.QST(GND),.B0Z(NET_902),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T25_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_20_padClk),.QRT(not_RESET_0_CAND2_BRSBL_20_tpGCLKBUF),.QST(GND),.T1I0(NET_62),.T1I1(m1_oper1_rdata_int[0]),.T1I2(NET_113_CAND4_BRSBL_20_tpGCLKBUF),.T1I3(m1_oper0_rdata_int[0]),.C1Z(NET_108),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_T25_2 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_20_padClk),.QRT(not_RESET_0_CAND2_BRSBL_20_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[0]),.T2I1(GND),.T2I2(nx11311z1_CAND5_BRSBL_20_tpGCLKBUF),.T2I3(m1_oper0_rdata_int[0]),.TB2S(GND),.Q2Z(tcdm_wdata_p2_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_T25_3 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_20_padClk),.QRT(not_RESET_0_CAND2_BRSBL_20_tpGCLKBUF),.QST(GND),.T3I0(nx11311z1_CAND5_BRSBL_20_tpGCLKBUF),.T3I1(GND),.T3I2(lint_WDATA_int[2]),.T3I3(m1_oper0_rdata_int[2]),.TB3S(GND),.Q3Z(tcdm_wdata_p2_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_T26_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B0I0(m1_oper0_rdata_int[6]),.B0I1(m1_oper1_rdata_int[6]),.B0I2(NET_113_CAND4_BRSBL_20_tpGCLKBUF),.B0I3(NET_62),.QCK(CLK_int_0__CAND0_BRSBL_20_padClk),.QRT(not_RESET_0_CAND2_BRSBL_20_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_rdata_int[12]),.T0I1(m1_oper0_rdata_int[12]),.T0I2(NET_113_CAND4_BRSBL_20_tpGCLKBUF),.T0I3(NET_62),.TB0S(GND),.B0Z(NET_800),.C0Z(NET_314),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_T26_1 (.tFragBitInfo(16'b0011001000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_20_padClk),.QRT(not_RESET_0_CAND2_BRSBL_20_tpGCLKBUF),.QST(GND),.T1I0(nx11311z1_CAND5_BRSBL_20_tpGCLKBUF),.T1I1(GND),.T1I2(m1_oper0_rdata_int[17]),.T1I3(lint_WDATA_int[17]),.TB1S(GND),.Q1Z(tcdm_wdata_p2_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_T26_2 (.tFragBitInfo(16'b0101010000000100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_20_padClk),.QRT(not_RESET_0_CAND2_BRSBL_20_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(m1_oper0_rdata_int[12]),.T2I2(nx11311z1_CAND5_BRSBL_20_tpGCLKBUF),.T2I3(lint_WDATA_int[12]),.TB2S(GND),.Q2Z(tcdm_wdata_p2_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_T26_3 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx30923z2),.QCK(CLK_int_0__CAND0_BRSBL_20_padClk),.QRT(not_RESET_0_CAND2_BRSBL_20_tpGCLKBUF),.QST(GND),.T3I0(m1_oper0_rdata_int[6]),.T3I1(lint_WDATA_int[6]),.T3I2(nx11311z1_CAND5_BRSBL_20_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p2_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_T30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_T30_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_T30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_T30_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m1_coef_rdata_int[17]),.T3I1(NET_111),.T3I2(m1_oper0_rdata_int[17]),.T3I3(NET_113_CAND4_BRSBL_20_tpGCLKBUF),.TB3S(GND),.C3Z(NET_454),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_U4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_112),.B0I1(m0_oper1_rdata_int[6]),.B0I2(NET_59_CAND5_TRSTL_21_tpGCLKBUF),.B0I3(m0_oper0_rdata_int[6]),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.B0Z(NET_801),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U4_2 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2_CAND3_TRSTL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.T2I0(nx11313z1_CAND2_TRSTL_21_tpGCLKBUF),.T2I1(m0_oper0_rdata_int[2]),.T2I2(lint_WDATA_int[2]),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_U4_3 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx41193z2_CAND3_TRSTL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[6]),.T3I1(GND),.T3I2(nx11313z1_CAND2_TRSTL_21_tpGCLKBUF),.T3I3(m0_oper0_rdata_int[6]),.TB3S(GND),.Q3Z(tcdm_wdata_p0_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_U5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_112),.B0I1(m0_oper1_rdata_int[2]),.B0I2(NET_59_CAND5_TRSTL_21_tpGCLKBUF),.B0I3(m0_oper0_rdata_int[2]),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.B0Z(NET_904),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U5_1 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx41193z2_CAND3_TRSTL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.T1I0(nx11313z1_CAND2_TRSTL_21_tpGCLKBUF),.T1I1(GND),.T1I2(lint_WDATA_int[12]),.T1I3(m0_oper0_rdata_int[12]),.TB1S(GND),.Q1Z(tcdm_wdata_p0_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_U5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_112),.B2I1(m0_oper1_rdata_int[12]),.B2I2(NET_59_CAND5_TRSTL_21_tpGCLKBUF),.B2I3(m0_oper0_rdata_int[12]),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.B2Z(NET_315),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_U6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U6_1 (.tFragBitInfo(16'b0000000010111000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx41193z2_CAND3_TRSTL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[17]),.T1I1(nx11313z1_CAND2_TRSTL_21_tpGCLKBUF),.T1I2(m0_oper0_rdata_int[17]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p0_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_U6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U6_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_U7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U7_1 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx41193z2_CAND3_TRSTL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.T1I0(m0_oper0_rdata_int[24]),.T1I1(nx11313z1_CAND2_TRSTL_21_tpGCLKBUF),.T1I2(lint_WDATA_int[24]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p0_dup_0[24]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_U7_2 (.tFragBitInfo(16'b0000111000000010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx41193z2_CAND3_TRSTL_21_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.T2I0(m0_oper0_rdata_int[26]),.T2I1(nx11313z1_CAND2_TRSTL_21_tpGCLKBUF),.T2I2(GND),.T2I3(lint_WDATA_int[26]),.TB2S(GND),.Q2Z(tcdm_wdata_p0_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_U7_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_21_padClk),.QRT(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_U10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(m0_oper1_wmode_dup_0[0]),.B0I1(fpgaio_in_int[6]),.B0I2(NET_143),.B0I3(NET_142),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B0Z(NET_810),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[14]),.Q1EN(nx41097z1),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_osel_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U10_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_143),.B2I1(fpgaio_in_int[7]),.B2I2(m0_oper1_wmode_dup_0[1]),.B2I3(NET_142),.CD2S(VCC),.Q2DI(lint_WDATA_int[9]),.Q2EN(nx41097z1),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T2I0(m1_m1_control[9]),.T2I1(NET_65),.T2I2(NET_37),.T2I3(tcdm_addr_p0_dup_0[9]),.TB2S(GND),.B2Z(NET_610),.C2Z(NET_251),.Q2Z(m1_m1_control[9]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_U10_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(tcdm_addr_p0_dup_0[14]),.T3I1(NET_65),.T3I2(NET_37),.T3I3(m1_m1_osel_dup_0),.C3Z(NET_360),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_U11_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T0I0(NET_37),.T0I1(tcdm_addr_p0_dup_0[10]),.T0I2(m1_m1_control[10]),.T0I3(NET_65),.TB0S(GND),.C0Z(NET_271),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[10]),.Q3EN(nx41097z1),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.Q3Z(m1_m1_control[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_U12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(m0_oper1_rdata_int[22]),.B0I1(m1_oper1_rdata_int[22]),.B0I2(NET_59),.B0I3(NET_62),.B0Z(NET_556),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U12_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(m0_m1_dataout_int[7]),.T1I1(NET_4),.T1I2(NET_116),.T1I3(NET_24),.C1Z(NET_611),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_U12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m0_oper0_rdata_int[17]),.B2I1(NET_112),.B2I2(NET_62),.B2I3(m1_oper1_rdata_int[17]),.B2Z(NET_455),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U12_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(m0_m1_dataout_int[6]),.T3I1(NET_4),.T3I2(NET_116),.T3I3(NET_24),.C3Z(NET_811),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_U13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0010000000000000),.B0I0(NET_610),.B0I1(GND),.B0I2(NET_608),.B0I3(NET_609),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.B0Z(NET_593),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx41097z1),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.Q1Z(m1_m1_mode_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_U13_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b1000000000000000),.B2I0(m0_m1_dataout_int[0]),.B2I1(NET_24),.B2I2(NET_4),.B2I3(NET_116),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T2I0(NET_37),.T2I1(NET_65),.T2I2(tcdm_addr_p0_dup_0[13]),.T2I3(m1_m1_mode_dup_0[1]),.TB2S(GND),.B2Z(NET_138),.C2Z(NET_348),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_U13_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(m0_m1_dataout_int[2]),.T3I1(NET_24),.T3I2(NET_4),.T3I3(NET_116),.C3Z(NET_913),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_U14_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[21]),.Q0EN(nx19726z1),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T0I0(NET_142),.T0I1(NET_140),.T0I2(m0_ram_control[22]),.T0I3(tcdm_result_p3[22]),.TB0S(GND),.C0Z(NET_557),.Q0Z(m0_ram_control[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U14_1 (.tFragBitInfo(16'b0000001100110011),.bFragBitInfo(16'b0000000000000111),.B1I0(NET_139),.B1I1(fpgaio_in_int[66]),.B1I2(tcdm_result_p3[2]),.B1I3(NET_913),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p3[2]),.T1I1(NET_913),.T1I2(NET_139),.T1I3(fpgaio_in_int[66]),.TB1S(NET_140),.C1Z(NET_911),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_U14_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0010000000000000),.B2I0(NET_810),.B2I1(GND),.B2I2(NET_808),.B2I3(NET_809),.CD2S(VCC),.Q2DI(lint_WDATA_int[22]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T2I0(NET_142),.T2I1(NET_140),.T2I2(tcdm_result_p3[21]),.T2I3(m0_ram_control[21]),.TB2S(GND),.B2Z(NET_793),.C2Z(NET_533),.Q2Z(m0_ram_control[22]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_U14_3 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_21_padClk),.QRT(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF),.QST(GND),.T3I0(NET_802),.T3I1(NET_800),.T3I2(GND),.T3I3(NET_801),.C3Z(NET_795),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_U15_0 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'b0000000000000000),.T0I0(NET_314),.T0I1(NET_315),.T0I2(NET_316),.T0I3(GND),.TB0S(GND),.C0Z(NET_309),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_U15_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_345),.T1I1(NET_348),.T1I2(NET_346),.T1I3(NET_347),.TB1S(GND),.C1Z(NET_349),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_U15_2 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0100000000000000),.B2I0(GND),.B2I1(NET_903),.B2I2(NET_904),.B2I3(NET_902),.T2I0(tcdm_result_p1[12]),.T2I1(NET_144),.T2I2(NET_145),.T2I3(m1_m1_dataout_int[12]),.TB2S(GND),.B2Z(NET_897),.C2Z(NET_322),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_U15_3 (.tFragBitInfo(16'b0001001100010011),.bFragBitInfo(16'b0000000000010011),.B3I0(NET_139),.B3I1(tcdm_result_p3[6]),.B3I2(fpgaio_in_int[70]),.B3I3(NET_811),.T3I0(fpgaio_in_int[70]),.T3I1(NET_811),.T3I2(NET_139),.T3I3(tcdm_result_p3[6]),.TB3S(NET_140),.C3Z(NET_809),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_U16_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_266),.B0I1(m1_m1_dataout_int[14]),.B0I2(tcdm_result_p1[14]),.B0I3(NET_42),.T0I0(NET_266),.T0I1(tcdm_addr_p1_dup_0[11]),.T0I2(NET_50),.T0I3(m1_m1_dataout_int[11]),.TB0S(GND),.B0Z(NET_370),.C0Z(NET_297),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_U16_1 (.tFragBitInfo(16'b0000001100110011),.bFragBitInfo(16'b0000000000000111),.B1I0(fpgaio_in_int[71]),.B1I1(NET_139),.B1I2(tcdm_result_p3[7]),.B1I3(NET_611),.T1I0(tcdm_result_p3[7]),.T1I1(NET_611),.T1I2(fpgaio_in_int[71]),.T1I3(NET_139),.TB1S(NET_140),.C1Z(NET_609),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_U16_2 (.tFragBitInfo(16'b0100010011001100),.bFragBitInfo(16'b0000010000001100),.B2I0(NET_69),.B2I1(NET_68),.B2I2(tcdm_addr_p3_dup_0[1]),.B2I3(m0_m1_dataout_int[1]),.T2I0(NET_69),.T2I1(NET_68),.T2I2(tcdm_addr_p3_dup_0[1]),.T2I3(m0_m1_dataout_int[1]),.TB2S(NET_70),.C2Z(NET_48),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_U16_3 (.tFragBitInfo(16'b0001000100110011),.bFragBitInfo(16'b0000000000010101),.B3I0(tcdm_result_p3[0]),.B3I1(NET_139),.B3I2(fpgaio_in_int[64]),.B3I3(NET_138),.T3I0(fpgaio_in_int[64]),.T3I1(NET_138),.T3I2(tcdm_result_p3[0]),.T3I3(NET_139),.TB3S(NET_140),.C3Z(NET_136),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_U17_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_1__CAND1_BRSTL_21_padClk),.QRT(not_RESET_1),.QST(GND),.T0I0(NET_249),.T0I1(NET_248),.T0I2(NET_251),.T0I3(NET_250),.TB0S(GND),.C0Z(NET_252),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U17_1 (.tFragBitInfo(16'b0000101010101010),.bFragBitInfo(16'b0000000001110000),.B1I0(cnt1[1]),.B1I1(NET_139),.B1I2(NET_453),.B1I3(tcdm_result_p3[17]),.QCK(CLK_int_1__CAND1_BRSTL_21_padClk),.QRT(not_RESET_1),.QST(GND),.T1I0(NET_453),.T1I1(tcdm_result_p3[17]),.T1I2(cnt1[1]),.T1I3(NET_139),.TB1S(NET_140),.C1Z(NET_449),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_U17_2 (.tFragBitInfo(16'b0000000100000010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(VCC),.QCK(CLK_int_1__CAND1_BRSTL_21_padClk),.QRT(not_RESET_1),.QST(GND),.T2I0(cnt1[1]),.T2I1(GND),.T2I2(GND),.T2I3(cnt1[0]),.TB2S(GND),.Q2Z(cnt1[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_U17_3 (.tFragBitInfo(16'b0001001000110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(VCC),.QCK(CLK_int_1__CAND1_BRSTL_21_padClk),.QRT(not_RESET_1),.QST(GND),.T3I0(cnt1[1]),.T3I1(GND),.T3I2(cnt1[2]),.T3I3(cnt1[0]),.TB3S(GND),.Q3Z(cnt1[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_U18_0 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0000000000000001),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(RESET_int[1]),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(GND),.QST(GND),.T0I0(fpgaio_out_dup_0[73]),.T0I1(NET_254),.T0I2(tcdm_addr_p3_dup_0[9]),.T0I3(NET_70),.TB0S(GND),.B0Z(not_RESET_1),.C0Z(NET_250),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U18_1 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(GND),.QST(GND),.T1I0(fpgaio_out_dup_0[69]),.T1I1(NET_254),.T1I2(GND),.T1I3(GND),.C1Z(NET_834),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_U18_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001001101011111),.B2I0(tcdm_addr_p3_dup_0[3]),.B2I1(NET_254),.B2I2(NET_70),.B2I3(fpgaio_out_dup_0[67]),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(GND),.QST(GND),.T2I0(fpgaio_out_dup_0[77]),.T2I1(NET_254),.T2I2(NET_70),.T2I3(tcdm_addr_p3_dup_0[13]),.TB2S(GND),.B2Z(NET_889),.C2Z(NET_346),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_U18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001000001010000),.B3I0(NET_834),.B3I1(tcdm_addr_p2_dup_0[5]),.B3I2(NET_835),.B3I3(NET_253),.CD3S(VCC),.Q3DI(lint_WDATA_int[31]),.Q3EN(nx40547z1),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(GND),.QST(GND),.T3I0(NET_835),.T3I1(NET_253),.T3I2(NET_834),.T3I3(tcdm_addr_p2_dup_0[5]),.TB3S(NET_836),.C3Z(NET_825),.Q3Z(tcdm_wen_p2_dup_0),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_U19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(lint_ADDR_int[4]),.B0I1(lint_ADDR_int[5]),.B0I2(lint_ADDR_int[6]),.B0I3(GND),.B0Z(NET_4),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U19_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_112),.T1I1(m1_oper1_rdata_int[24]),.T1I2(NET_62_CAND3_BRSTL_21_tpGCLKBUF),.T1I3(m0_oper0_rdata_int[24]),.C1Z(NET_624),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_U19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_112),.B2I1(m1_oper1_rdata_int[26]),.B2I2(NET_62_CAND3_BRSTL_21_tpGCLKBUF),.B2I3(m0_oper0_rdata_int[26]),.B2Z(NET_663),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_U23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND2_BRSTL_21_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U23_1 (.tFragBitInfo(16'b0000001100000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1EN(VCC),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND2_BRSTL_21_tpGCLKBUF),.QST(GND),.T1I0(nx50994z1),.T1I1(GND),.T1I2(GND),.T1I3(nx50994z2),.TB1S(GND),.Q1Z(launch_p3),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.Q1DI(GND),.T1CO());

	LOGIC_2 QL_INST_U23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000001110000),.B2I0(p3_fsm[0]),.B2I1(launch_p3),.B2I2(control_in_int[3]),.B2I3(last_control[3]),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND2_BRSTL_21_tpGCLKBUF),.QST(GND),.B2Z(nx50994z1),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(control_in_int[3]),.Q3EN(VCC),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(not_RESET_0_CAND2_BRSTL_21_tpGCLKBUF),.QST(GND),.Q3Z(last_control[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_U24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100110100001100),.B0I0(p3_cnt[0]),.B0I1(control_in_int[17]),.B0I2(p3_cnt[1]),.B0I3(control_in_int[16]),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(GND),.QST(GND),.B0Z(NET_158),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_U24_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(GND),.QST(GND),.T1I0(NET_152),.T1I1(NET_151),.T1I2(NET_150),.T1I3(GND),.C1Z(NET_148),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_U24_2 (.tFragBitInfo(16'b0000000100000010),.bFragBitInfo(16'b1000001001000001),.B2I0(p3_cnt[0]),.B2I1(control_in_int[17]),.B2I2(p3_cnt[1]),.B2I3(control_in_int[16]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(GND),.QST(GND),.T2I0(p3_cnt[1]),.T2I1(GND),.T2I2(p3_fsm[0]),.T2I3(p3_cnt[0]),.TB2S(GND),.B2Z(NET_150),.Q2Z(p3_cnt[1]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_U24_3 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSTL_21_padClk),.QRT(GND),.QST(GND),.T3I0(GND),.T3I1(GND),.T3I2(p3_fsm[0]),.T3I3(p3_cnt[0]),.TB3S(GND),.Q3Z(p3_cnt[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_U25_0 (.tFragBitInfo(16'b0000000001101100),.bFragBitInfo(16'b1000001001000001),.B0I0(control_in_int[19]),.B0I1(p3_cnt[2]),.B0I2(control_in_int[18]),.B0I3(p3_cnt[3]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSBL_21_padClk),.QRT(GND),.QST(GND),.T0I0(p3_cnt[1]),.T0I1(p3_cnt[2]),.T0I2(p3_cnt[0]),.T0I3(p3_fsm_0__CAND1_BRSBL_21_tpGCLKBUF),.TB0S(GND),.B0Z(NET_152),.Q0Z(p3_cnt[2]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U25_1 (.tFragBitInfo(16'b0001001100000001),.bFragBitInfo(16'b0100110111111111),.B1I0(control_in_int[18]),.B1I1(p3_cnt[2]),.B1I2(NET_158),.B1I3(control_in_int[19]),.QCK(CLK_int_0__CAND0_BRSBL_21_padClk),.QRT(GND),.QST(GND),.T1I0(NET_158),.T1I1(control_in_int[19]),.T1I2(control_in_int[18]),.T1I3(p3_cnt[2]),.TB1S(p3_cnt[3]),.C1Z(NET_157),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_U25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(p3_cnt[1]),.B2I1(p3_cnt[2]),.B2I2(p3_cnt[0]),.B2I3(p3_cnt[3]),.QCK(CLK_int_0__CAND0_BRSBL_21_padClk),.QRT(GND),.QST(GND),.B2Z(NET_740),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_U25_3 (.tFragBitInfo(16'b0011001100000000),.bFragBitInfo(16'b0000000001101100),.B3I0(p3_cnt[0]),.B3I1(p3_cnt[3]),.B3I2(p3_cnt[1]),.B3I3(p3_fsm_0__CAND1_BRSBL_21_tpGCLKBUF),.CD3S(GND),.Q3DI(GND),.Q3EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSBL_21_padClk),.QRT(GND),.QST(GND),.T3I0(p3_cnt[1]),.T3I1(p3_fsm_0__CAND1_BRSBL_21_tpGCLKBUF),.T3I2(p3_cnt[0]),.T3I3(p3_cnt[3]),.TB3S(p3_cnt[2]),.Q3Z(p3_cnt[3]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_U27_0 (.tFragBitInfo(16'b0000000100000100),.bFragBitInfo(16'b0000000000000001),.B0I0(p3_cnt[9]),.B0I1(p3_cnt[8]),.B0I2(p3_cnt[10]),.B0I3(p3_cnt[11]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSBL_21_padClk),.QRT(GND),.QST(GND),.T0I0(GND),.T0I1(NET_739),.T0I2(p3_fsm_0__CAND1_BRSBL_21_tpGCLKBUF),.T0I3(p3_cnt[8]),.TB0S(GND),.B0Z(NET_155),.Q0Z(p3_cnt[8]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_U27_1 (.tFragBitInfo(16'b0000000000010010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSBL_21_padClk),.QRT(GND),.QST(GND),.T1I0(NET_819),.T1I1(p3_fsm_0__CAND1_BRSBL_21_tpGCLKBUF),.T1I2(p3_cnt[10]),.T1I3(GND),.TB1S(GND),.Q1Z(p3_cnt[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_U27_2 (.tFragBitInfo(16'b0000011000001010),.bFragBitInfo(16'b0000100000000000),.B2I0(p3_cnt[9]),.B2I1(NET_739),.B2I2(GND),.B2I3(p3_cnt[8]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSBL_21_padClk),.QRT(GND),.QST(GND),.T2I0(p3_cnt[9]),.T2I1(NET_739),.T2I2(p3_fsm_0__CAND1_BRSBL_21_tpGCLKBUF),.T2I3(p3_cnt[8]),.TB2S(GND),.B2Z(NET_819),.Q2Z(p3_cnt[9]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_U27_3 (.tFragBitInfo(16'b0001001100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSBL_21_padClk),.QRT(GND),.QST(GND),.T3I0(NET_819),.T3I1(p3_fsm_0__CAND1_BRSBL_21_tpGCLKBUF),.T3I2(p3_cnt[10]),.T3I3(p3_cnt[11]),.TB3S(GND),.Q3Z(p3_cnt[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_V8_0 (.tFragBitInfo(16'b0000010100000100),.bFragBitInfo(16'b0000011100000000),.B0I0(p1_fsm_0__CAND4_TRSTL_22_tpGCLKBUF),.B0I1(launch_p1),.B0I2(last_control[1]),.B0I3(control_in_int[1]),.CD0S(GND),.Q0EN(VCC),.QCK(CLK_int_0__CAND0_TRSTL_22_padClk),.QRT(not_RESET_0_CAND1_TRSTL_22_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(nx50996z2),.T0I2(GND),.T0I3(nx50996z1),.TB0S(GND),.B0Z(nx50996z1),.Q0Z(launch_p1),.B0CO(),.C0Z(),.Q0DI(GND),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_V8_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_22_padClk),.QRT(not_RESET_0_CAND1_TRSTL_22_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(control_in_int[1]),.Q2EN(VCC),.QCK(CLK_int_0__CAND0_TRSTL_22_padClk),.QRT(not_RESET_0_CAND1_TRSTL_22_tpGCLKBUF),.QST(GND),.Q2Z(last_control[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V8_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_22_padClk),.QRT(not_RESET_0_CAND1_TRSTL_22_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx19726z1),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.Q2Z(m0_oper1_wmode_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[7]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.Q3Z(m0_oper1_wmode_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[20]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p1[20]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V12_0 (.tFragBitInfo(16'b0001000101010101),.bFragBitInfo(16'b0000000100000101),.B0I0(NET_505),.B0I1(NET_145),.B0I2(m0_ram_control[19]),.B0I3(tcdm_result_p1[19]),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T0I0(NET_505),.T0I1(NET_145),.T0I2(m0_ram_control[19]),.T0I3(tcdm_result_p1[19]),.TB0S(NET_142),.C0Z(NET_496),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_V12_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[19]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p1_dup_0[17]),.T1I1(NET_116),.T1I2(NET_35),.T1I3(NET_4),.C1Z(NET_458),.Q1Z(m0_ram_control[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_V12_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000100000000),.B2I0(lint_ADDR_int[3]),.B2I1(GND),.B2I2(lint_ADDR_int[11]),.B2I3(lint_ADDR_int[2]),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T2I0(NET_4),.T2I1(NET_116),.T2I2(NET_35),.T2I3(tcdm_addr_p1_dup_0[19]),.TB2S(GND),.B2Z(NET_116),.C2Z(NET_505),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_V12_3 (.tFragBitInfo(16'b0001000100110011),.bFragBitInfo(16'b0000000000010101),.B3I0(m0_ram_control[17]),.B3I1(tcdm_result_p1[17]),.B3I2(NET_145),.B3I3(NET_458),.CD3S(VCC),.Q3DI(lint_WDATA_int[17]),.Q3EN(nx19726z1),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T3I0(NET_145),.T3I1(NET_458),.T3I2(m0_ram_control[17]),.T3I3(tcdm_result_p1[17]),.TB3S(NET_142),.C3Z(NET_448),.Q3Z(m0_ram_control[17]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_V13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100000000000000),.B0I0(GND),.B0I1(NET_35),.B0I2(NET_4),.B0I3(NET_116),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B0Z(NET_115),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[22]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p1[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V13_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T3I0(NET_145),.T3I1(NET_144),.T3I2(m1_m1_dataout_int[7]),.T3I3(tcdm_result_p1[7]),.C3Z(NET_608),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_V14_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_145),.B0I1(tcdm_result_p1[18]),.B0I2(NET_142),.B0I3(m0_ram_control[18]),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T0I0(NET_468),.T0I1(NET_467),.T0I2(NET_469),.T0I3(NET_470),.TB0S(GND),.B0Z(NET_469),.C0Z(NET_471),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_V14_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[18]),.Q1EN(nx19726z1),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T1I0(tcdm_result_p1[2]),.T1I1(NET_144),.T1I2(m1_m1_dataout_int[2]),.T1I3(NET_145),.C1Z(NET_910),.Q1Z(m0_ram_control[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_V14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0100110001011111),.B2I0(fpgaio_in_int[18]),.B2I1(NET_472),.B2I2(NET_143),.B2I3(NET_473),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B2Z(NET_468),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V14_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T3I0(tcdm_result_p1[6]),.T3I1(NET_144),.T3I2(NET_145),.T3I3(m1_m1_dataout_int[6]),.C3Z(NET_808),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_V15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[27]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p1[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V15_1 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(lint_ADDR_int[11]),.T1I2(NET_53),.T1I3(NET_35),.TB1S(GND),.C1Z(NET_473),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_V15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(m1_m1_dataout_int[0]),.B2I1(NET_144),.B2I2(NET_145),.B2I3(tcdm_result_p1[0]),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B2Z(NET_135),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_42),.B0I1(NET_51),.B0I2(tcdm_result_p1[9]),.B0I3(i_events[9]),.CD0S(VCC),.Q0DI(lint_WDATA_int[9]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B0Z(NET_232),.Q0Z(i_events[9]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V16_1 (.tFragBitInfo(16'b0011111100000000),.bFragBitInfo(16'b0000010000001100),.B1I0(m0_m1_dataout_int[4]),.B1I1(NET_867),.B1I2(tcdm_addr_p2_dup_0[4]),.B1I3(NET_69),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p2_dup_0[4]),.T1I1(NET_69),.T1I2(m0_m1_dataout_int[4]),.T1I3(NET_867),.TB1S(NET_253),.C1Z(NET_863),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_V16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_42),.B2I1(tcdm_result_p1[13]),.B2I2(NET_253),.B2I3(tcdm_addr_p2_dup_0[13]),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.B2Z(NET_331),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V16_3 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_22_padClk),.QRT(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_33),.T3I2(NET_53),.T3I3(GND),.C3Z(NET_253),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_V17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V17_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.T2I0(tcdm_result_p3[18]),.T2I1(NET_139),.T2I2(cnt1[2]),.T2I3(NET_140),.TB2S(GND),.C2Z(NET_467),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_V17_3 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_29),.T3I1(NET_53),.T3I2(GND),.T3I3(GND),.C3Z(NET_70),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_V18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_253),.B0I1(tcdm_addr_p2_dup_0[15]),.B0I2(NET_254),.B0I3(fpgaio_out_dup_0[79]),.B0Z(NET_408),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V18_2 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_40),.T2I1(GND),.T2I2(GND),.T2I3(NET_29),.TB2S(GND),.C2Z(NET_51),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_V18_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(NET_407),.T3I1(NET_408),.T3I2(NET_406),.T3I3(GND),.C3Z(NET_395),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_V19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V19_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[3]),.T1I1(NET_4),.T1I2(NET_35),.T1I3(tcdm_be_p3_dup_0[0]),.C1Z(NET_526),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_V19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[16]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[4]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p3[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[23]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p3[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[0]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p3[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_V23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[12]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V24_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[14]),.T1I1(NET_198),.T1I2(NET_10),.T1I3(GND),.C1Z(nx3850z2),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_V24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V24_3 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[30]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_22_padClk),.QRT(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[14]),.T3I1(NET_198),.T3I2(GND),.T3I3(NET_79),.TB3S(GND),.C3Z(NET_508),.Q3Z(tcdm_result_p3[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_V25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V25_1 (.tFragBitInfo(16'b1000000000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_153),.T1I1(NET_154),.T1I2(control_in_int[20]),.T1I3(p3_cnt[4]),.C1Z(NET_151),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_V25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_V25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_V26_0 (.tFragBitInfo(16'b0000011000001100),.bFragBitInfo(16'b0000001000000000),.B0I0(p3_cnt[4]),.B0I1(GND),.B0I2(GND),.B0I3(p3_cnt[5]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSBL_22_padClk),.QRT(GND),.QST(GND),.T0I0(p3_cnt[4]),.T0I1(p3_cnt[5]),.T0I2(p3_fsm_0__CAND1_BRSBL_22_tpGCLKBUF),.T0I3(NET_740),.TB0S(GND),.B0Z(NET_741),.Q0Z(p3_cnt[5]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_V26_1 (.tFragBitInfo(16'b1101111101010101),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_22_padClk),.QRT(GND),.QST(GND),.T1I0(NET_155),.T1I1(NET_160),.T1I2(NET_154),.T1I3(NET_159),.C1Z(NET_156),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_V26_2 (.tFragBitInfo(16'b0000000100000010),.bFragBitInfo(16'b1011111100001011),.B2I0(p3_cnt[4]),.B2I1(control_in_int[20]),.B2I2(control_in_int[21]),.B2I3(p3_cnt[5]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSBL_22_padClk),.QRT(GND),.QST(GND),.T2I0(p3_cnt[4]),.T2I1(p3_fsm_0__CAND1_BRSBL_22_tpGCLKBUF),.T2I2(GND),.T2I3(NET_740),.TB2S(GND),.B2Z(NET_160),.Q2Z(p3_cnt[4]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_V26_3 (.tFragBitInfo(16'b0000000010000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_22_padClk),.QRT(GND),.QST(GND),.T3I0(NET_155),.T3I1(p3_cnt[5]),.T3I2(control_in_int[21]),.T3I3(GND),.C3Z(NET_153),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_V27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_741),.B0I1(NET_740),.B0I2(p3_cnt[6]),.B0I3(p3_cnt[7]),.QCK(CLK_int_0__CAND0_BRSBL_22_padClk),.QRT(GND),.QST(GND),.B0Z(NET_739),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_V27_1 (.tFragBitInfo(16'b1111011100110001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_22_padClk),.QRT(GND),.QST(GND),.T1I0(control_in_int[22]),.T1I1(control_in_int[23]),.T1I2(p3_cnt[6]),.T1I3(p3_cnt[7]),.C1Z(NET_159),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_V27_2 (.tFragBitInfo(16'b0001001000110000),.bFragBitInfo(16'b1000010000100001),.B2I0(control_in_int[22]),.B2I1(control_in_int[23]),.B2I2(p3_cnt[6]),.B2I3(p3_cnt[7]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSBL_22_padClk),.QRT(GND),.QST(GND),.T2I0(NET_741),.T2I1(p3_fsm_0__CAND1_BRSBL_22_tpGCLKBUF),.T2I2(p3_cnt[6]),.T2I3(NET_740),.TB2S(GND),.B2Z(NET_154),.Q2Z(p3_cnt[6]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_V27_3 (.tFragBitInfo(16'b0011001100000000),.bFragBitInfo(16'b0000000001101100),.B3I0(NET_740),.B3I1(p3_cnt[7]),.B3I2(NET_741),.B3I3(p3_fsm_0__CAND1_BRSBL_22_tpGCLKBUF),.CD3S(GND),.Q3DI(GND),.Q3EN(nx56739z2),.QCK(CLK_int_0__CAND0_BRSBL_22_padClk),.QRT(GND),.QST(GND),.T3I0(NET_741),.T3I1(p3_fsm_0__CAND1_BRSBL_22_tpGCLKBUF),.T3I2(NET_740),.T3I3(p3_cnt[7]),.TB3S(p3_cnt[6]),.Q3Z(p3_cnt[7]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_W2_0 (.tFragBitInfo(16'b0000011000001100),.bFragBitInfo(16'b0000000010000000),.B0I0(NET_219),.B0I1(p1_cnt[9]),.B0I2(p1_cnt[8]),.B0I3(GND),.CD0S(GND),.Q0DI(GND),.Q0EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.T0I0(NET_219),.T0I1(p1_cnt[9]),.T0I2(p1_fsm_0__CAND4_TRSTL_23_tpGCLKBUF),.T0I3(p1_cnt[8]),.TB0S(GND),.B0Z(NET_548),.Q0Z(p1_cnt[9]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W2_1 (.tFragBitInfo(16'b0000000100010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.T1I0(p1_fsm_0__CAND4_TRSTL_23_tpGCLKBUF),.T1I1(GND),.T1I2(NET_548),.T1I3(p1_cnt[10]),.TB1S(GND),.Q1Z(p1_cnt[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_W2_2 (.tFragBitInfo(16'b0001010001000100),.bFragBitInfo(16'b0000000000000001),.B2I0(p1_cnt[9]),.B2I1(p1_cnt[11]),.B2I2(p1_cnt[8]),.B2I3(p1_cnt[10]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.T2I0(p1_fsm_0__CAND4_TRSTL_23_tpGCLKBUF),.T2I1(p1_cnt[11]),.T2I2(NET_548),.T2I3(p1_cnt[10]),.TB2S(GND),.B2Z(NET_185),.Q2Z(p1_cnt[11]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_W2_3 (.tFragBitInfo(16'b0000000000010010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.T3I0(NET_219),.T3I1(p1_fsm_0__CAND4_TRSTL_23_tpGCLKBUF),.T3I2(p1_cnt[8]),.T3I3(GND),.TB3S(GND),.Q3Z(p1_cnt[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_W3_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W3_2 (.tFragBitInfo(16'b0101000001010000),.bFragBitInfo(16'b0001010001010000),.B2I0(p1_fsm_0__CAND4_TRSTL_23_tpGCLKBUF),.B2I1(p1_cnt[0]),.B2I2(p1_cnt[3]),.B2I3(p1_cnt[1]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.T2I0(p1_fsm_0__CAND4_TRSTL_23_tpGCLKBUF),.T2I1(p1_cnt[0]),.T2I2(p1_cnt[3]),.T2I3(p1_cnt[1]),.TB2S(p1_cnt[2]),.Q2Z(p1_cnt[3]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_W3_3 (.tFragBitInfo(16'b0000000010110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.T3I0(control_in_int[23]),.T3I1(p1_cnt[7]),.T3I2(NET_185),.T3I3(GND),.C3Z(NET_176),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_W4_0 (.tFragBitInfo(16'b0000000100000100),.bFragBitInfo(16'b0000101100001010),.B0I0(control_in_int[17]),.B0I1(p1_cnt[0]),.B0I2(p1_cnt[1]),.B0I3(control_in_int[16]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.T0I0(GND),.T0I1(p1_cnt[0]),.T0I2(p1_fsm_0__CAND4_TRSTL_23_tpGCLKBUF),.T0I3(p1_cnt[1]),.TB0S(GND),.B0Z(NET_184),.Q0Z(p1_cnt[1]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W4_1 (.tFragBitInfo(16'b0000000000000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.T1I0(p1_cnt[3]),.T1I1(control_in_int[19]),.T1I2(GND),.T1I3(GND),.C1Z(NET_182),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_W4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000001000000000),.B2I0(control_in_int[17]),.B2I1(p1_cnt[0]),.B2I2(GND),.B2I3(control_in_int[16]),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.B2Z(NET_183),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W4_3 (.tFragBitInfo(16'b0000111100000001),.bFragBitInfo(16'b0000000000000100),.B3I0(NET_182),.B3I1(p1_cnt[2]),.B3I2(NET_183),.B3I3(NET_184),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(GND),.T3I0(NET_183),.T3I1(NET_184),.T3I2(NET_182),.T3I3(p1_cnt[2]),.TB3S(control_in_int[18]),.C3Z(NET_181),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_W5_0 (.tFragBitInfo(16'b0000000000001010),.bFragBitInfo(16'b0000000000101111),.B0I0(NET_176),.B0I1(NET_175),.B0I2(p1_fsm[2]),.B0I3(p1_fsm[1]),.CD0S(GND),.Q0EN(nx3668z1),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.T0I0(p1_fsm_0__CAND4_TRSTL_23_tpGCLKBUF),.T0I1(GND),.T0I2(tcdm_wen_p1_dup_0),.T0I3(GND),.TB0S(GND),.B0Z(NET_174),.Q0Z(p1_fsm[1]),.B0CO(),.C0Z(),.Q0DI(GND),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W5_2 (.tFragBitInfo(16'b0001000100010000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2EN(nx3668z1),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(GND),.T2I2(nx1674z1),.T2I3(p1_fsm[1]),.TB2S(GND),.Q2Z(p1_fsm[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.Q2DI(GND),.T2CO());

	LOGIC_3 QL_INST_W5_3 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.T3I0(NET_176),.T3I1(NET_175),.T3I2(tcdm_wen_p1_dup_0),.T3I3(p1_fsm[4]),.TB3S(GND),.C3Z(nx1674z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_W6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W6_1 (.tFragBitInfo(16'b0000000000001110),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1EN(nx3668z1),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.T1I0(nx11312z5),.T1I1(nx3668z8),.T1I2(GND),.T1I3(GND),.TB1S(GND),.Q1Z(p1_fsm[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.Q1DI(GND),.T1CO());

	LOGIC_2 QL_INST_W6_2 (.tFragBitInfo(16'b0000101100000000),.bFragBitInfo(16'b0000000010110000),.B2I0(NET_175),.B2I1(NET_176),.B2I2(p1_fsm[2]),.B2I3(GND),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.T2I0(NET_175),.T2I1(NET_176),.T2I2(GND),.T2I3(p1_fsm[4]),.TB2S(GND),.B2Z(nx11312z5),.C2Z(nx3668z8),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_W6_3 (.tFragBitInfo(16'b0000000011111000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(GND),.QST(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.T3I0(tcdm_req_p0_dup_0),.T3I1(p0_fsm[4]),.T3I2(nx45272z2),.T3I3(GND),.C3Z(nx42281z2),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_W7_0 (.tFragBitInfo(16'b0100010001010000),.bFragBitInfo(16'b0110101010101010),.B0I0(tcdm_addr_p0_dup_0[17]),.B0I1(tcdm_addr_p0_dup_0[15]),.B0I2(tcdm_addr_p0_dup_0[16]),.B0I3(NET_736),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(lint_WDATA_int[17]),.T0I2(NET_742),.T0I3(nx45272z2),.TB0S(GND),.B0Z(NET_742),.Q0Z(tcdm_addr_p0_dup_0[17]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W7_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p0_dup_0[17]),.T1I1(tcdm_addr_p0_dup_0[15]),.T1I2(tcdm_addr_p0_dup_0[16]),.T1I3(NET_736),.C1Z(NET_735),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_W7_2 (.tFragBitInfo(16'b1011000111100100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.T2I0(nx45272z2),.T2I1(tcdm_addr_p0_dup_0[18]),.T2I2(lint_WDATA_int[18]),.T2I3(NET_735),.TB2S(GND),.Q2Z(tcdm_addr_p0_dup_0[18]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_W7_3 (.tFragBitInfo(16'b0100010000000101),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTL_23_padClk),.QRT(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(lint_WDATA_int[2]),.T3I2(tcdm_addr_p0_dup_0[2]),.T3I3(nx45272z2),.TB3S(GND),.Q3Z(tcdm_addr_p0_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_W9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W9_2 (.tFragBitInfo(16'b0000011000001010),.bFragBitInfo(16'b1111011011111010),.B2I0(tcdm_addr_p0_dup_0[4]),.B2I1(tcdm_addr_p0_dup_0[2]),.B2I2(nx45272z2),.B2I3(tcdm_addr_p0_dup_0[3]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p0_dup_0[4]),.T2I1(tcdm_addr_p0_dup_0[2]),.T2I2(nx45272z2),.T2I3(tcdm_addr_p0_dup_0[3]),.TB2S(lint_WDATA_int[4]),.Q2Z(tcdm_addr_p0_dup_0[4]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_W9_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_W10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[3]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p1[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[1]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p1[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_W11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[5]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p1[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[8]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p1[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx45272z2),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p0_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_W12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[17]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p1[17]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[19]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p1[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_W13_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(GND),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[31]),.Q1EN(nx40545z1),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_wen_p0_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(fpgaio_in_int[50]),.B2I1(NET_115),.B2I2(NET_114),.B2I3(tcdm_addr_p1_dup_0[18]),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(GND),.QST(GND),.B2Z(NET_470),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W13_3 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(GND),.QST(GND),.T3I0(NET_90),.T3I1(NET_81),.T3I2(NET_91),.T3I3(GND),.TB3S(GND),.C3Z(nx45272z2),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_W14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_900),.B1I1(NET_897),.B1I2(NET_899),.B1I3(NET_898),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.T1I0(NET_899),.T1I1(NET_898),.T1I2(NET_900),.T1I3(NET_897),.TB1S(NET_901),.C1Z(NET_893),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_W14_2 (.tFragBitInfo(16'b0000110111011101),.bFragBitInfo(16'b0000011101110111),.B2I0(NET_107),.B2I1(tcdm_addr_p0_dup_0[2]),.B2I2(NET_106),.B2I3(tcdm_result_p2[2]),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[9]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.T2I0(NET_107),.T2I1(tcdm_be_p0_dup_0[3]),.T2I2(NET_106),.T2I3(tcdm_result_p2[23]),.TB2S(GND),.B2Z(NET_899),.C2Z(NET_587),.Q2Z(tcdm_result_p1[9]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_W14_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[30]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.T3I0(NET_115),.T3I1(NET_114),.T3I2(tcdm_addr_p1_dup_0[2]),.T3I3(fpgaio_in_int[34]),.C3Z(NET_900),.Q3Z(tcdm_result_p1[30]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_W15_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_140),.B0I1(tcdm_result_p3[26]),.B0I2(tcdm_result_p1[26]),.B0I3(NET_145),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.T0I0(NET_50),.T0I1(NET_51),.T0I2(tcdm_addr_p1_dup_0[15]),.T0I3(i_events[15]),.TB0S(GND),.B0Z(NET_665),.C0Z(NET_407),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W15_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[15]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.T1I0(NET_140),.T1I1(tcdm_result_p1[28]),.T1I2(tcdm_result_p3[28]),.T1I3(NET_145),.C1Z(NET_707),.Q1Z(i_events[15]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_W15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(tcdm_result_p3[29]),.B2I1(tcdm_result_p1[29]),.B2I2(NET_140),.B2I3(NET_145),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[28]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.B2Z(NET_730),.Q2Z(tcdm_result_p1[28]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W15_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[26]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.T3I0(NET_140),.T3I1(tcdm_result_p1[24]),.T3I2(tcdm_result_p3[24]),.T3I3(NET_145),.C3Z(NET_626),.Q3Z(tcdm_result_p1[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_W16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx60509z1),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.Q0Z(i_events[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W16_1 (.tFragBitInfo(16'b0101000011110000),.bFragBitInfo(16'b0000000000101010),.B1I0(NET_49),.B1I1(tcdm_addr_p1_dup_0[1]),.B1I2(NET_50),.B1I3(i_events[1]),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.T1I0(NET_50),.T1I1(i_events[1]),.T1I2(NET_49),.T1I3(tcdm_addr_p1_dup_0[1]),.TB1S(NET_51),.C1Z(NET_45),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_W16_2 (.tFragBitInfo(16'b0100110001001100),.bFragBitInfo(16'b0000000001001100),.B2I0(fpgaio_out_dup_0[68]),.B2I1(NET_927),.B2I2(NET_254),.B2I3(tcdm_addr_p1_dup_0[4]),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.T2I0(fpgaio_out_dup_0[68]),.T2I1(NET_927),.T2I2(NET_254),.T2I3(tcdm_addr_p1_dup_0[4]),.TB2S(NET_50),.C2Z(NET_928),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_W16_3 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_23_padClk),.QRT(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[4]),.T3I1(lint_ADDR_int[6]),.T3I2(lint_ADDR_int[5]),.T3I3(lint_ADDR_int[3]),.TB3S(GND),.C3Z(NET_53),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_W17_0 (.tFragBitInfo(16'b0001000000000000),.bFragBitInfo(16'b0000000000100000),.B0I0(NET_29),.B0I1(GND),.B0I2(NET_40),.B0I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[5]),.T0I1(lint_ADDR_int[4]),.T0I2(lint_ADDR_int[3]),.T0I3(lint_ADDR_int[6]),.TB0S(GND),.B0Z(NET_105),.C0Z(NET_52),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W17_1 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[23]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(NET_33),.T1I2(NET_53),.T1I3(lint_ADDR_int[11]),.TB1S(GND),.C1Z(NET_104),.Q1Z(tcdm_result_p2[23]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_W17_2 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'b0000000000001000),.B2I0(NET_52),.B2I1(NET_33),.B2I2(GND),.B2I3(lint_ADDR_int[11]),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(NET_33),.T2I2(GND),.T2I3(NET_52),.TB2S(GND),.B2Z(NET_118),.C2Z(NET_254),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_W17_3 (.tFragBitInfo(16'b0111011111111111),.bFragBitInfo(16'b0001111101011111),.B3I0(NET_53),.B3I1(NET_52),.B3I2(NET_33),.B3I3(fpgaio_out_dup_0[65]),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[2]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.T3I0(NET_33),.T3I1(fpgaio_out_dup_0[65]),.T3I2(NET_53),.T3I3(NET_52),.TB3S(tcdm_addr_p2_dup_0[1]),.C3Z(NET_49),.Q3Z(tcdm_result_p2[2]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_W18_0 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0001010100111111),.B0I0(NET_119),.B0I1(fpgaio_out_dup_0[66]),.B0I2(NET_118),.B0I3(tcdm_addr_p3_dup_0[2]),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.T0I0(NET_53),.T0I1(NET_29),.T0I2(GND),.T0I3(tcdm_addr_p3_dup_0[14]),.TB0S(GND),.B0Z(NET_901),.C0Z(NET_363),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W18_1 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.T1I0(NET_53),.T1I1(NET_29),.T1I2(GND),.T1I3(tcdm_addr_p3_dup_0[11]),.TB1S(GND),.C1Z(NET_290),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_W18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000001000),.B2I0(NET_53),.B2I1(NET_29),.B2I2(lint_ADDR_int[11]),.B2I3(GND),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.B2Z(NET_119),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W18_3 (.tFragBitInfo(16'b0011111111111111),.bFragBitInfo(16'b0000011111111111),.B3I0(NET_40),.B3I1(i_events[4]),.B3I2(tcdm_addr_p3_dup_0[4]),.B3I3(NET_29),.CD3S(VCC),.Q3DI(lint_WDATA_int[4]),.Q3EN(nx60509z1),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.T3I0(tcdm_addr_p3_dup_0[4]),.T3I1(NET_29),.T3I2(NET_40),.T3I3(i_events[4]),.TB3S(NET_53),.C3Z(NET_927),.Q3Z(i_events[4]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_W20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[29]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p3[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_W21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[22]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p3[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[6]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p3[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[25]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[25]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_W22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[9]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p3[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[21]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p3[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[31]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_W23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000001),.B0I0(GND),.B0I1(p3_fsm[0]),.B0I2(GND),.B0I3(GND),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[18]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.B0Z(not_p3_fsm_0),.Q0Z(tcdm_result_p3[18]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W23_1 (.tFragBitInfo(16'b0000000000110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1EN(nx20469z1),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(not_p3_fsm_0),.T1I2(tcdm_wen_p3_dup_0),.T1I3(GND),.TB1S(GND),.Q1Z(p3_fsm[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.Q1DI(GND),.T1CO());

	LOGIC_2 QL_INST_W23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W23_3 (.tFragBitInfo(16'b0000000000001100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3EN(nx20469z1),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(p3_fsm[0]),.T3I2(tcdm_wen_p3_dup_0),.T3I3(GND),.TB3S(GND),.Q3Z(p3_fsm[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.Q3DI(GND),.T3CO());

	LOGIC_0 QL_INST_W24_0 (.tFragBitInfo(16'b0010000011110000),.bFragBitInfo(16'b0010000010100000),.B0I0(tcdm_gnt_p3_int),.B0I1(NET_149),.B0I2(NET_818),.B0I3(p3_fsm[2]),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.T0I0(tcdm_gnt_p3_int),.T0I1(NET_149),.T0I2(NET_818),.T0I3(p3_fsm[2]),.TB0S(p3_fsm[3]),.C0Z(nx56739z2),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W24_1 (.tFragBitInfo(16'b0000010100000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1EN(nx20469z1),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.T1I0(GND),.T1I1(p3_fsm[2]),.T1I2(GND),.T1I3(p3_fsm[4]),.TB1S(GND),.Q1Z(p3_fsm[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.Q1DI(GND),.T1CO());

	LOGIC_2 QL_INST_W24_2 (.tFragBitInfo(16'b0000110100001111),.bFragBitInfo(16'b0000000000010000),.B2I0(GND),.B2I1(p3_fsm[1]),.B2I2(RESET_int[0]),.B2I3(p3_fsm[4]),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.T2I0(launch_p3),.T2I1(p3_fsm[2]),.T2I2(NET_508),.T2I3(p3_fsm[0]),.TB2S(GND),.B2Z(NET_818),.C2Z(NET_509),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_W24_3 (.tFragBitInfo(16'b0000000100000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_23_padClk),.QRT(GND),.QST(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF),.T3I0(launch_p3),.T3I1(GND),.T3I2(GND),.T3I3(p3_fsm[0]),.C3Z(NET_221),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_W25_0 (.tFragBitInfo(16'b0000000011001000),.bFragBitInfo(16'b0000110000000100),.B0I0(NET_151),.B0I1(NET_156),.B0I2(GND),.B0I3(NET_157),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T0I0(NET_220),.T0I1(tcdm_valid_p3_int),.T0I2(p3_fsm[3]),.T0I3(GND),.TB0S(GND),.B0Z(NET_149),.C0Z(nx30664z1),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(p3_fsm[1]),.Q1EN(nx20469z1),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.Q1Z(p3_fsm[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W25_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000010001),.B2I0(NET_220),.B2I1(NET_221),.B2I2(p3_fsm[3]),.B2I3(NET_222),.CD2S(VCC),.Q2DI(p3_fsm[3]),.Q2EN(nx20469z1),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T2I0(NET_220),.T2I1(NET_221),.T2I2(p3_fsm[3]),.T2I3(NET_222),.TB2S(NET_148),.C2Z(nx20469z1),.Q2Z(p3_fsm[4]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_W25_3 (.tFragBitInfo(16'b0011000010110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T3I0(NET_151),.T3I1(NET_156),.T3I2(p3_fsm[2]),.T3I3(NET_157),.TB3S(GND),.C3Z(NET_222),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_W26_0 (.tFragBitInfo(16'b0000000000000010),.bFragBitInfo(16'b1100110011011100),.B0I0(p3_fsm[1]),.B0I1(nx3850z2_CAND3_BRSBL_23_tpGCLKBUF),.B0I2(NET_926),.B0I3(p3_fsm[2]),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T0I0(p3_fsm[4]),.T0I1(GND),.T0I2(NET_223),.T0I3(GND),.TB0S(GND),.B0Z(nx64401z2),.C0Z(NET_220),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W26_1 (.tFragBitInfo(16'b0000000000001110),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1EN(VCC),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T1I0(nx30664z1),.T1I1(nx3850z2_CAND3_BRSBL_23_tpGCLKBUF),.T1I2(GND),.T1I3(GND),.TB1S(GND),.Q1Z(m1_oper1_we_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.Q1DI(GND),.T1CO());

	LOGIC_2 QL_INST_W26_2 (.tFragBitInfo(16'b1101111111001110),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T2I0(p3_fsm[4]),.T2I1(nx3850z2_CAND3_BRSBL_23_tpGCLKBUF),.T2I2(NET_223),.T2I3(p3_fsm[3]),.TB2S(GND),.C2Z(nx3786z2),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_W26_3 (.tFragBitInfo(16'b0011000000110001),.bFragBitInfo(16'b0000000000001011),.B3I0(m1_oper1_we_dup_0),.B3I1(p3_fsm[3]),.B3I2(p3_fsm[4]),.B3I3(NET_221),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T3I0(p3_fsm[4]),.T3I1(NET_221),.T3I2(m1_oper1_we_dup_0),.T3I3(p3_fsm[3]),.TB3S(NET_223),.C3Z(NET_926),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_W27_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W27_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W27_2 (.tFragBitInfo(16'b1000001000000000),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_225),.T2I1(m1_oper1_waddr_dup_0[0]),.T2I2(control_in_int[14]),.T2I3(NET_224),.TB2S(GND),.C2Z(NET_223),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_W27_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_W28_0 (.tFragBitInfo(16'b1100110100000001),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_waddr_dup_0[2]),.T0I1(nx3850z2_CAND3_BRSBL_23_tpGCLKBUF),.T0I2(p3_fsm_0__CAND1_BRSBL_23_tpGCLKBUF),.T0I3(lint_ADDR_int[2]),.TB0S(GND),.Q0Z(m1_oper1_waddr_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_W28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_W28_2 (.tFragBitInfo(16'b1000001001000001),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_waddr_dup_0[2]),.T2I1(control_in_int[17]),.T2I2(m1_oper1_waddr_dup_0[3]),.T2I3(control_in_int[16]),.TB2S(GND),.C2Z(NET_225),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_W28_3 (.tFragBitInfo(16'b1000001001000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T3I0(m1_oper1_waddr_dup_0[1]),.T3I1(control_in_int[18]),.T3I2(m1_oper1_waddr_dup_0[4]),.T3I3(control_in_int[15]),.TB3S(GND),.C3Z(NET_228),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_W30_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_W30_1 (.tFragBitInfo(16'b1010000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[4]),.T1I1(NET_891),.T1I2(nx3850z2_CAND3_BRSBL_23_tpGCLKBUF),.T1I3(p3_fsm_0__CAND1_BRSBL_23_tpGCLKBUF),.TB1S(GND),.Q1Z(m1_oper1_waddr_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_W30_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010101000000),.B2I0(GND),.B2I1(m1_oper1_waddr_dup_0[3]),.B2I2(m1_oper1_waddr_dup_0[2]),.B2I3(m1_oper1_waddr_dup_0[4]),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.B2Z(NET_891),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_W30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_23_padClk),.QRT(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X1_0 (.tFragBitInfo(16'b1101100010001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T0I0(NET_77),.T0I1(lint_ADDR_int[7]),.T0I2(p1_fsm[4]),.T0I3(p1_cnt[5]),.TB0S(GND),.Q0Z(m0_oper1_raddr_dup_0[7]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X1_1 (.tFragBitInfo(16'b1100110010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T1I0(p1_fsm[3]),.T1I1(lint_ADDR_int[7]),.T1I2(p1_cnt[5]),.T1I3(nx25587z2),.TB1S(GND),.Q1Z(m0_oper1_waddr_dup_0[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_X1_2 (.tFragBitInfo(16'b1110101001000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T2I0(NET_77),.T2I1(p1_cnt[2]),.T2I2(p1_fsm[4]),.T2I3(lint_ADDR_int[4]),.TB2S(GND),.Q2Z(m0_oper1_raddr_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_X1_3 (.tFragBitInfo(16'b1111100000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T3I0(p1_fsm[3]),.T3I1(p1_cnt[2]),.T3I2(nx25587z2),.T3I3(lint_ADDR_int[4]),.TB3S(GND),.Q3Z(m0_oper1_waddr_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_X2_0 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_214),.B0I1(NET_212),.B0I2(p1_cnt[6]),.B0I3(p1_cnt[7]),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T0I0(p1_cnt[4]),.T0I1(GND),.T0I2(GND),.T0I3(p1_cnt[5]),.TB0S(GND),.B0Z(NET_219),.C0Z(NET_214),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X2_1 (.tFragBitInfo(16'b0000111100000000),.bFragBitInfo(16'b0001010001000100),.B1I0(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.B1I1(p1_cnt[7]),.B1I2(NET_214),.B1I3(NET_212),.CD1S(GND),.Q1DI(GND),.Q1EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T1I0(NET_214),.T1I1(NET_212),.T1I2(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.T1I3(p1_cnt[7]),.TB1S(p1_cnt[6]),.Q1Z(p1_cnt[7]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_X2_2 (.tFragBitInfo(16'b0000000000000110),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T2I0(p1_cnt[4]),.T2I1(NET_212),.T2I2(GND),.T2I3(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.TB2S(GND),.Q2Z(p1_cnt[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_X2_3 (.tFragBitInfo(16'b0000000001111000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T3I0(NET_214),.T3I1(NET_212),.T3I2(p1_cnt[6]),.T3I3(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.TB3S(GND),.Q3Z(p1_cnt[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_X3_0 (.tFragBitInfo(16'b0000011000001010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T0I0(p1_cnt[5]),.T0I1(p1_cnt[4]),.T0I2(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.T0I3(NET_212),.TB0S(GND),.Q0Z(p1_cnt[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X3_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T1I0(p1_cnt[1]),.T1I1(p1_cnt[3]),.T1I2(p1_cnt[2]),.T1I3(p1_cnt[0]),.TB1S(GND),.C1Z(NET_212),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_X3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X3_3 (.tFragBitInfo(16'b1010111100100011),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T3I0(p1_cnt[7]),.T3I1(control_in_int[22]),.T3I2(control_in_int[23]),.T3I3(p1_cnt[6]),.C3Z(NET_177),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_X4_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b1011000010111011),.B0I0(p1_cnt[5]),.B0I1(control_in_int[21]),.B0I2(p1_cnt[4]),.B0I3(control_in_int[20]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T0I0(GND),.T0I1(p1_cnt[0]),.T0I2(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.T0I3(GND),.TB0S(GND),.B0Z(NET_179),.Q0Z(p1_cnt[0]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X4_1 (.tFragBitInfo(16'b0010101000001010),.bFragBitInfo(16'b1101000011010000),.B1I0(NET_178),.B1I1(NET_179),.B1I2(NET_177),.B1I3(NET_180),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T1I0(NET_177),.T1I1(NET_180),.T1I2(NET_178),.T1I3(NET_179),.TB1S(NET_181),.C1Z(NET_175),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_X4_2 (.tFragBitInfo(16'b0000011000001010),.bFragBitInfo(16'b1111010100110001),.B2I0(p1_cnt[4]),.B2I1(p1_cnt[3]),.B2I2(control_in_int[20]),.B2I3(control_in_int[19]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx14855z2),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T2I0(p1_cnt[2]),.T2I1(p1_cnt[0]),.T2I2(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.T2I3(p1_cnt[1]),.TB2S(GND),.B2Z(NET_180),.Q2Z(p1_cnt[2]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_X4_3 (.tFragBitInfo(16'b1100010011110101),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(GND),.QST(GND),.T3I0(p1_cnt[6]),.T3I1(control_in_int[21]),.T3I2(control_in_int[22]),.T3I3(p1_cnt[5]),.C3Z(NET_178),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_X5_0 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'b0000000000001000),.B0I0(RESET_int[0]),.B0I1(NET_174),.B0I2(p1_fsm[4]),.B0I3(NET_213),.T0I0(lint_ADDR_int[12]),.T0I1(NET_78),.T0I2(NET_79),.T0I3(GND),.TB0S(GND),.B0Z(nx14855z2),.C0Z(NET_77),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO());

	LOGIC_1 QL_INST_X5_1 (.tFragBitInfo(16'b1111010011110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(lint_ADDR_int[12]),.T1I1(NET_78),.T1I2(p1_fsm[3]),.T1I3(NET_10),.TB1S(GND),.C1Z(nx39177z2),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO());

	LOGIC_2 QL_INST_X5_2 (.tFragBitInfo(16'b1010111010101010),.bFragBitInfo(16'b0000000000000001),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(tcdm_wen_p1_dup_0),.T2I0(NET_481),.T2I1(NET_78),.T2I2(lint_ADDR_int[12]),.T2I3(NET_10),.TB2S(GND),.B2Z(not_tcdm_wen_p1),.C2Z(nx35588z2),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_X5_3 (.tFragBitInfo(16'b1111111101000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T3I0(lint_ADDR_int[12]),.T3I1(NET_78),.T3I2(NET_79),.T3I3(NET_215),.TB3S(GND),.C3Z(nx18281z3),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO());

	LOGIC_0 QL_INST_X6_0 (.tFragBitInfo(16'b0001000100010000),.bFragBitInfo(16'b1010110000100000),.B0I0(m0_oper1_we_dup_0),.B0I1(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.B0I2(p1_fsm[3]),.B0I3(launch_p1),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T0I0(tcdm_gnt_p1_int),.T0I1(GND),.T0I2(p1_fsm[3]),.T0I3(p1_fsm[2]),.TB0S(GND),.B0Z(NET_481),.C0Z(NET_213),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X6_1 (.tFragBitInfo(16'b0100010001001100),.bFragBitInfo(16'b0011111100000000),.B1I0(NET_176),.B1I1(p1_fsm[3]),.B1I2(NET_213),.B1I3(NET_507),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T1I0(NET_213),.T1I1(NET_507),.T1I2(NET_176),.T1I3(p1_fsm[3]),.TB1S(NET_175),.C1Z(nx3668z1),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_X6_2 (.tFragBitInfo(16'b0011000010111000),.bFragBitInfo(16'b1100110011101100),.B2I0(p1_fsm[4]),.B2I1(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.B2I2(NET_176),.B2I3(NET_175),.CD2S(GND),.Q2DI(GND),.Q2EN(nx3668z1),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T2I0(NET_176),.T2I1(p1_fsm[2]),.T2I2(p1_fsm[3]),.T2I3(NET_175),.TB2S(GND),.B2Z(nx677z1),.C2Z(nx65216z1),.Q2Z(p1_fsm[4]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_X6_3 (.tFragBitInfo(16'b0000000000001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3EN(nx3668z1),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T3I0(nx677z1),.T3I1(GND),.T3I2(not_tcdm_wen_p1),.T3I3(GND),.TB3S(GND),.Q3Z(p1_fsm[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.Q3DI(GND),.T3CO());

	LOGIC_0 QL_INST_X7_0 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b0000100000000000),.B0I0(tcdm_wen_p1_dup_0),.B0I1(p1_fsm[4]),.B0I2(GND),.B0I3(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T0I0(NET_10),.T0I1(NET_78),.T0I2(lint_ADDR_int[12]),.T0I3(GND),.TB0S(GND),.B0Z(nx25587z1),.C0Z(nx25587z2),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X7_1 (.tFragBitInfo(16'b1010111100100011),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T1I0(launch_p1),.T1I1(p1_fsm[4]),.T1I2(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.T1I3(tcdm_valid_p1_int),.C1Z(NET_507),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_X7_2 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T2I0(nx25587z2),.T2I1(lint_WDATA_int[31]),.T2I2(GND),.T2I3(tcdm_rdata_p1_int[31]),.TB2S(GND),.Q2Z(m0_oper1_wdata_dup_0[31]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_X7_3 (.tFragBitInfo(16'b0000000000110010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3EN(VCC),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T3I0(nx25587z2),.T3I1(GND),.T3I2(nx25587z1),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper1_we_dup_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.Q3DI(GND),.T3CO());

	LOGIC_0 QL_INST_X8_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1110001001000000),.B0I0(p1_fsm[4]),.B0I1(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.B0I2(launch_p1),.B0I3(tcdm_req_p1_dup_0),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.B0Z(NET_215),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X8_1 (.tFragBitInfo(16'b0000000000001110),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1EN(nx11312z3),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T1I0(nx11312z1),.T1I1(nx65216z1),.T1I2(GND),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_req_p1_dup_0),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.Q1DI(GND),.T1CO());

	LOGIC_2 QL_INST_X8_2 (.tFragBitInfo(16'b0011001000010000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T2I0(nx25587z2),.T2I1(GND),.T2I2(tcdm_rdata_p1_int[30]),.T2I3(lint_WDATA_int[30]),.TB2S(GND),.Q2Z(m0_oper1_wdata_dup_0[30]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_X8_3 (.tFragBitInfo(16'b1111111110111010),.bFragBitInfo(16'b1111000011111010),.B3I0(tcdm_gnt_p1_int),.B3I1(NET_174),.B3I2(nx11312z1),.B3I3(tcdm_fmo_p1_int),.QCK(CLK_int_0__CAND0_TRSTL_24_padClk),.QRT(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF),.QST(GND),.T3I0(nx11312z1),.T3I1(tcdm_fmo_p1_int),.T3I2(tcdm_gnt_p1_int),.T3I3(NET_174),.TB3S(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF),.C3Z(nx11312z3),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_X10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[10]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p1[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[7]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p1[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[11]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p1[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[12]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p1[12]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X11_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X11_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[15]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p1[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[21]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p1[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[6]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p1[6]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X13_0 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[24]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.T0I0(RESET_int[0]),.T0I1(GND),.T0I2(GND),.T0I3(nx45272z2),.TB0S(GND),.C0Z(nx40545z1),.Q0Z(tcdm_result_p1[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X13_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[31]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p1[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X13_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[23]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.T2I0(NET_90),.T2I1(NET_91),.T2I2(GND),.T2I3(lint_ADDR_int[2]),.TB2S(GND),.C2Z(NET_89),.Q2Z(tcdm_result_p1[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_X13_3 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.T3I0(NET_90),.T3I1(NET_91),.T3I2(GND),.T3I3(lint_ADDR_int[2]),.C3Z(nx12973z2),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_X14_0 (.tFragBitInfo(16'b1101000011011101),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_90),.B0I1(NET_91),.B0I2(lint_ADDR_int[2]),.B0I3(RESET_int[0]),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(GND),.QST(GND),.T0I0(NET_115),.T0I1(tcdm_be_p1_dup_0[1]),.T0I2(tcdm_be_p3_dup_0[1]),.T0I3(NET_473),.TB0S(GND),.B0Z(nx40546z1),.C0Z(NET_539),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X14_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(GND),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X14_2 (.tFragBitInfo(16'b1101000011011101),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[31]),.Q2EN(nx40546z1),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(GND),.QST(GND),.T2I0(NET_115),.T2I1(tcdm_be_p1_dup_0[3]),.T2I2(tcdm_be_p3_dup_0[3]),.T2I3(NET_473),.TB2S(GND),.C2Z(NET_581),.Q2Z(tcdm_wen_p1_dup_0),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_X14_3 (.tFragBitInfo(16'b1100010011110101),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(GND),.QST(GND),.T3I0(NET_115),.T3I1(tcdm_be_p3_dup_0[2]),.T3I2(tcdm_be_p1_dup_0[2]),.T3I3(NET_473),.TB3S(GND),.C3Z(NET_562),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_X15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_99),.B1I1(NET_101),.B1I2(NET_100),.B1I3(NET_102),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[13]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.T1I0(NET_100),.T1I1(NET_102),.T1I2(NET_99),.T1I3(NET_101),.TB1S(NET_103),.C1Z(NET_95),.Q1Z(tcdm_result_p1[13]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_X15_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(fpgaio_in_int[32]),.B2I1(tcdm_addr_p1_dup_0[0]),.B2I2(NET_114),.B2I3(NET_115),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[29]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.B2Z(NET_102),.Q2Z(tcdm_result_p1[29]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X15_3 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[25]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBL_24_padClk),.QRT(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF),.QST(GND),.T3I0(NET_106),.T3I1(NET_107),.T3I2(tcdm_result_p2[0]),.T3I3(tcdm_addr_p0_dup_0[0]),.C3Z(NET_101),.Q3Z(tcdm_result_p1[25]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_X16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001000000000000),.B2I0(GND),.B2I1(GND),.B2I2(lint_ADDR_int[7]),.B2I3(NET_10),.B2Z(NET_3),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[0]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p2[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X17_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.T1I0(NET_104),.T1I1(NET_105),.T1I2(tcdm_addr_p2_dup_0[0]),.T1I3(i_events[0]),.C1Z(NET_100),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_X17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[0]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q2Z(i_events[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(tcdm_addr_p3_dup_0[0]),.B0I1(fpgaio_out_dup_0[64]),.B0I2(NET_119),.B0I3(NET_118),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B0Z(NET_103),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X18_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[12]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p2[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_90),.B2I1(NET_10),.B2I2(NET_1),.B2I3(NET_2),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B2Z(nx40548z2),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[0]),.Q3EN(nx40548z2),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_addr_p3_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[14]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p3[14]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[17]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[17]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[10]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p3[10]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X21_0 (.tFragBitInfo(16'b0000100000001101),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60936z2),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.T0I0(nx40548z2),.T0I1(lint_WDATA_int[2]),.T0I2(GND),.T0I3(tcdm_addr_p3_dup_0[2]),.TB0S(GND),.Q0Z(tcdm_addr_p3_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[1]),.Q1EN(nx40548z2),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_addr_p3_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[11]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p3[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X22_0 (.tFragBitInfo(16'b1100110011111111),.bFragBitInfo(16'b0100110001011111),.B0I0(NET_1),.B0I1(tcdm_fmo_p3_int),.B0I2(NET_2),.B0I3(tcdm_gnt_p3_int),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[28]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.T0I0(NET_1),.T0I1(tcdm_fmo_p3_int),.T0I2(NET_2),.T0I3(tcdm_gnt_p3_int),.TB0S(NET_3),.C0Z(NET_161),.Q0Z(tcdm_result_p3[28]),.B0CO(),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X22_1 (.tFragBitInfo(16'b0001010001010000),.bFragBitInfo(16'b1111011011111010),.B1I0(tcdm_addr_p3_dup_0[4]),.B1I1(tcdm_addr_p3_dup_0[3]),.B1I2(nx40548z2),.B1I3(tcdm_addr_p3_dup_0[2]),.CD1S(GND),.Q1DI(GND),.Q1EN(nx60936z2),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.T1I0(nx40548z2),.T1I1(tcdm_addr_p3_dup_0[2]),.T1I2(tcdm_addr_p3_dup_0[4]),.T1I3(tcdm_addr_p3_dup_0[3]),.TB1S(lint_WDATA_int[4]),.Q1Z(tcdm_addr_p3_dup_0[4]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_X22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[1]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[1]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X22_3 (.tFragBitInfo(16'b0100000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_3),.T3I2(NET_2),.T3I3(NET_1),.C3Z(NET_0),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_X23_0 (.tFragBitInfo(16'b1111111100010000),.bFragBitInfo(16'b1111111100010101),.B0I0(NET_148),.B0I1(NET_149),.B0I2(p3_fsm[2]),.B0I3(NET_0),.CD0S(GND),.Q0DI(GND),.Q0EN(nx11310z3),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.T0I0(NET_148),.T0I1(NET_149),.T0I2(p3_fsm[2]),.T0I3(NET_0),.TB0S(p3_fsm[3]),.Q0Z(tcdm_req_p3_dup_0),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X23_1 (.tFragBitInfo(16'b1111111100100000),.bFragBitInfo(16'b1100111011101110),.B1I0(tcdm_gnt_p3_int),.B1I1(nx40548z2),.B1I2(p3_fsm[2]),.B1I3(NET_149),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[27]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.T1I0(p3_fsm[2]),.T1I1(NET_149),.T1I2(tcdm_gnt_p3_int),.T1I3(nx40548z2),.TB1S(p3_fsm[3]),.C1Z(nx60936z2),.Q1Z(tcdm_result_p3[27]),.B1CO(),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_X23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X23_3 (.tFragBitInfo(16'b0001111100001111),.bFragBitInfo(16'b0101011101011111),.B3I0(NET_161),.B3I1(p3_fsm[2]),.B3I2(NET_148),.B3I3(NET_149),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[7]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.T3I0(NET_148),.T3I1(NET_149),.T3I2(NET_161),.T3I3(p3_fsm[2]),.TB3S(p3_fsm[3]),.C3Z(nx11310z3),.Q3Z(tcdm_result_p3[7]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_X24_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[5]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p3[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_X24_1 (.tFragBitInfo(16'b0000000001110011),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.T1I0(NET_149),.T1I1(NET_509),.T1I2(NET_510),.T1I3(GND),.C1Z(nx36808z2),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_X24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X24_3 (.tFragBitInfo(16'b0000000001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[19]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTL_24_padClk),.QRT(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF),.QST(GND),.T3I0(tcdm_fmo_p3_int),.T3I1(p3_fsm[2]),.T3I2(tcdm_gnt_p3_int),.T3I3(NET_221),.TB3S(GND),.C3Z(NET_510),.Q3Z(tcdm_result_p3[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_X26_0 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T0I0(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.T0I1(lint_WDATA_int[31]),.T0I2(GND),.T0I3(tcdm_rdata_p3_int[31]),.TB0S(GND),.Q0Z(m1_oper1_wdata_dup_0[31]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X26_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p3_int[21]),.T1I1(lint_WDATA_int[21]),.T1I2(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(m1_oper1_wdata_dup_0[21]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_X26_2 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T2I0(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.T2I1(GND),.T2I2(lint_WDATA_int[29]),.T2I3(tcdm_rdata_p3_int[29]),.TB2S(GND),.Q2Z(m1_oper1_wdata_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_X26_3 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p3_int[19]),.T3I1(lint_WDATA_int[19]),.T3I2(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper1_wdata_dup_0[19]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_X27_0 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000010),.B0I0(m1_oper1_waddr_dup_0[1]),.B0I1(GND),.B0I2(GND),.B0I3(p3_fsm_0__CAND1_BRSBL_24_tpGCLKBUF),.CD0S(GND),.Q0EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(nx16644z1),.T0I2(nx16644z2),.T0I3(lint_ADDR_int[1]),.TB0S(GND),.B0Z(nx16644z1),.Q0Z(m1_oper1_waddr_dup_0[1]),.B0CO(),.C0Z(),.Q0DI(GND),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X27_1 (.tFragBitInfo(16'b0000000000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(p3_fsm_0__CAND1_BRSBL_24_tpGCLKBUF),.T1I2(m1_oper1_waddr_dup_0[0]),.T1I3(GND),.TB1S(GND),.C1Z(nx17641z1),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_X27_2 (.tFragBitInfo(16'b0100010001010000),.bFragBitInfo(16'b0000000000000001),.B2I0(GND),.B2I1(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.B2I2(GND),.B2I3(GND),.CD2S(GND),.Q2DI(GND),.Q2EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_WDATA_int[25]),.T2I2(tcdm_rdata_p3_int[25]),.T2I3(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.TB2S(GND),.B2Z(nx16644z2),.Q2Z(m1_oper1_wdata_dup_0[25]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_X27_3 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[0]),.T3I1(nx16644z2),.T3I2(nx17641z1),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper1_waddr_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.Q3DI(GND),.T3CO());

	LOGIC_0 QL_INST_X28_0 (.tFragBitInfo(16'b1000001001000001),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_waddr_dup_0[7]),.T0I1(control_in_int[23]),.T0I2(m1_oper1_waddr_dup_0[9]),.T0I3(control_in_int[21]),.TB0S(GND),.C0Z(NET_229),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X28_1 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[30]),.T1I1(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.T1I2(GND),.T1I3(tcdm_rdata_p3_int[30]),.TB1S(GND),.Q1Z(m1_oper1_wdata_dup_0[30]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_X28_2 (.tFragBitInfo(16'b1000010000100001),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_227),.B2I1(NET_229),.B2I2(NET_226),.B2I3(NET_228),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T2I0(control_in_int[19]),.T2I1(control_in_int[20]),.T2I2(m1_oper1_waddr_dup_0[5]),.T2I3(m1_oper1_waddr_dup_0[6]),.TB2S(GND),.B2Z(NET_224),.C2Z(NET_227),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_X28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X29_0 (.tFragBitInfo(16'b1010000010101100),.bFragBitInfo(16'b0000011000001010),.B0I0(m1_oper1_waddr_dup_0[7]),.B0I1(NET_303),.B0I2(GND),.B0I3(m1_oper1_waddr_dup_0[6]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[7]),.T0I1(NET_529),.T0I2(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.T0I3(p3_fsm_0__CAND1_BRSBL_24_tpGCLKBUF),.TB0S(GND),.B0Z(NET_529),.Q0Z(m1_oper1_waddr_dup_0[7]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X29_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X29_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X29_3 (.tFragBitInfo(16'b1010000010101100),.bFragBitInfo(16'b1010000010110001),.B3I0(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.B3I1(p3_fsm_0__CAND1_BRSBL_24_tpGCLKBUF),.B3I2(lint_ADDR_int[6]),.B3I3(NET_303),.CD3S(GND),.Q3DI(GND),.Q3EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T3I0(lint_ADDR_int[6]),.T3I1(NET_303),.T3I2(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.T3I3(p3_fsm_0__CAND1_BRSBL_24_tpGCLKBUF),.TB3S(m1_oper1_waddr_dup_0[6]),.Q3Z(m1_oper1_waddr_dup_0[6]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_X30_0 (.tFragBitInfo(16'b1000101110001000),.bFragBitInfo(16'b1000100010001011),.B0I0(lint_ADDR_int[3]),.B0I1(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.B0I2(p3_fsm_0__CAND1_BRSBL_24_tpGCLKBUF),.B0I3(m1_oper1_waddr_dup_0[2]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[3]),.T0I1(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.T0I2(p3_fsm_0__CAND1_BRSBL_24_tpGCLKBUF),.T0I3(m1_oper1_waddr_dup_0[2]),.TB0S(m1_oper1_waddr_dup_0[3]),.Q0Z(m1_oper1_waddr_dup_0[3]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X30_1 (.tFragBitInfo(16'b1100111000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T1I0(NET_218),.T1I1(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF),.T1I2(p3_fsm_0__CAND1_BRSBL_24_tpGCLKBUF),.T1I3(lint_ADDR_int[5]),.TB1S(GND),.Q1Z(m1_oper1_waddr_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_X30_2 (.tFragBitInfo(16'b0111100011110000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_waddr_dup_0[3]),.T2I1(m1_oper1_waddr_dup_0[4]),.T2I2(m1_oper1_waddr_dup_0[5]),.T2I3(m1_oper1_waddr_dup_0[2]),.TB2S(GND),.C2Z(NET_218),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_X30_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_X31_0 (.tFragBitInfo(16'b1010110010100000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx36808z2),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.T0I0(lint_ADDR_int[4]),.T0I1(p3_fsm[2]),.T0I2(NET_508),.T0I3(NET_530),.TB0S(GND),.Q0Z(m1_oper1_raddr_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_X31_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_X31_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_X31_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBL_24_padClk),.QRT(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y1_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y1_1 (.tFragBitInfo(16'b1110010010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T1I0(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF),.T1I1(p1_cnt[8]),.T1I2(lint_ADDR_int[10]),.T1I3(p1_fsm[3]),.TB1S(GND),.Q1Z(m0_oper1_waddr_dup_0[10]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y1_2 (.tFragBitInfo(16'b1111000010001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T2I0(p1_fsm[4]),.T2I1(p1_cnt[8]),.T2I2(lint_ADDR_int[10]),.T2I3(NET_77),.TB2S(GND),.Q2Z(m0_oper1_raddr_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y1_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y2_0 (.tFragBitInfo(16'b1101100010001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T0I0(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF),.T0I1(lint_ADDR_int[11]),.T0I2(p1_fsm[3]),.T0I3(p1_cnt[9]),.TB0S(GND),.Q0Z(m0_oper1_waddr_dup_0[11]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y2_1 (.tFragBitInfo(16'b1101100010001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T1I0(NET_77),.T1I1(lint_ADDR_int[11]),.T1I2(p1_fsm[4]),.T1I3(p1_cnt[9]),.TB1S(GND),.Q1Z(m0_oper1_raddr_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y2_2 (.tFragBitInfo(16'b1110110000100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T2I0(p1_fsm[4]),.T2I1(NET_77),.T2I2(p1_cnt[7]),.T2I3(lint_ADDR_int[9]),.TB2S(GND),.Q2Z(m0_oper1_raddr_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y2_3 (.tFragBitInfo(16'b1110110000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T3I0(p1_cnt[7]),.T3I1(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF),.T3I2(p1_fsm[3]),.T3I3(lint_ADDR_int[9]),.TB3S(GND),.Q3Z(m0_oper1_waddr_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y3_0 (.tFragBitInfo(16'b1101100010001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T0I0(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF),.T0I1(lint_ADDR_int[3]),.T0I2(p1_cnt[1]),.T0I3(p1_fsm[3]),.TB0S(GND),.Q0Z(m0_oper1_waddr_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y3_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y3_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y3_3 (.tFragBitInfo(16'b1110101001000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T3I0(NET_77),.T3I1(p1_fsm[4]),.T3I2(p1_cnt[1]),.T3I3(lint_ADDR_int[3]),.TB3S(GND),.Q3Z(m0_oper1_raddr_dup_0[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y4_3 (.tFragBitInfo(16'b0000110000001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36058z2_CAND4_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T3I0(m0_oper1_rdata_int[28]),.T3I1(lint_WDATA_int[28]),.T3I2(GND),.T3I3(nx11312z1_CAND3_TRSTR_25_tpGCLKBUF),.TB3S(GND),.Q3Z(tcdm_wdata_p1_dup_0[28]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y5_0 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx39177z2_CAND5_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p1_int[24]),.T0I1(GND),.T0I2(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF),.T0I3(lint_WDATA_int[24]),.TB0S(GND),.Q0Z(m0_oper1_wdata_dup_0[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y5_2 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx36058z2_CAND4_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[29]),.T2I1(nx11312z1_CAND3_TRSTR_25_tpGCLKBUF),.T2I2(GND),.T2I3(m0_oper1_rdata_int[29]),.TB2S(GND),.Q2Z(tcdm_wdata_p1_dup_0[29]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y5_3 (.tFragBitInfo(16'b0000000001010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(p1_fsm[2]),.T3I2(nx11312z1_CAND3_TRSTR_25_tpGCLKBUF),.T3I3(GND),.C3Z(nx36058z2),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_Y6_0 (.tFragBitInfo(16'b0000111000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx36058z2_CAND4_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T0I0(m0_oper1_rdata_int[23]),.T0I1(nx11312z1_CAND3_TRSTR_25_tpGCLKBUF),.T0I2(GND),.T0I3(lint_WDATA_int[23]),.TB0S(GND),.Q0Z(tcdm_wdata_p1_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y6_1 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx39177z2_CAND5_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T1I0(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF),.T1I1(GND),.T1I2(lint_WDATA_int[26]),.T1I3(tcdm_rdata_p1_int[26]),.TB1S(GND),.Q1Z(m0_oper1_wdata_dup_0[26]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y6_2 (.tFragBitInfo(16'b0000111000000100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx39177z2_CAND5_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T2I0(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF),.T2I1(tcdm_rdata_p1_int[23]),.T2I2(GND),.T2I3(lint_WDATA_int[23]),.TB2S(GND),.Q2Z(m0_oper1_wdata_dup_0[23]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y6_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx39177z2_CAND5_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[22]),.T3I1(tcdm_rdata_p1_int[22]),.T3I2(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper1_wdata_dup_0[22]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y7_0 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'b0010000000000000),.B0I0(tcdm_addr_p0_dup_0[12]),.B0I1(GND),.B0I2(tcdm_addr_p0_dup_0[13]),.B0I3(tcdm_addr_p0_dup_0[14]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx36058z2_CAND4_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[30]),.T0I1(GND),.T0I2(nx11312z1_CAND3_TRSTR_25_tpGCLKBUF),.T0I3(m0_oper1_rdata_int[30]),.TB0S(GND),.B0Z(NET_738),.Q0Z(tcdm_wdata_p1_dup_0[30]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(tcdm_addr_p0_dup_0[10]),.B1I1(tcdm_addr_p0_dup_0[11]),.B1I2(NET_737),.B1I3(NET_738),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T1I0(NET_737),.T1I1(NET_738),.T1I2(tcdm_addr_p0_dup_0[10]),.T1I3(tcdm_addr_p0_dup_0[11]),.TB1S(tcdm_addr_p0_dup_0[9]),.C1Z(NET_736),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_Y7_2 (.tFragBitInfo(16'b1100110001011010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p0_dup_0[15]),.T2I1(lint_WDATA_int[15]),.T2I2(NET_736),.T2I3(nx45272z2),.TB2S(GND),.Q2Z(tcdm_addr_p0_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y7_3 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36058z2_CAND4_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T3I0(nx11312z1_CAND3_TRSTR_25_tpGCLKBUF),.T3I1(lint_WDATA_int[31]),.T3I2(m0_oper1_rdata_int[31]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p1_dup_0[31]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y8_0 (.tFragBitInfo(16'b1100010111001010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T0I0(tcdm_addr_p0_dup_0[2]),.T0I1(lint_WDATA_int[3]),.T0I2(nx45272z2),.T0I3(tcdm_addr_p0_dup_0[3]),.TB0S(GND),.Q0Z(tcdm_addr_p0_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y8_1 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx39177z2_CAND5_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p1_int[19]),.T1I1(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF),.T1I2(lint_WDATA_int[19]),.T1I3(GND),.TB1S(GND),.Q1Z(m0_oper1_wdata_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y8_3 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx39177z2_CAND5_TRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_25_padClk),.QRT(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p1_int[20]),.T3I1(lint_WDATA_int[20]),.T3I2(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper1_wdata_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y9_0 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[29]),.T0I1(tcdm_rdata_p1_int[29]),.T0I2(nx25587z2),.T0I3(GND),.TB0S(GND),.Q0Z(m0_oper1_wdata_dup_0[29]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y9_1 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[25]),.T1I1(GND),.T1I2(nx25587z2),.T1I3(tcdm_rdata_p1_int[25]),.TB1S(GND),.Q1Z(m0_oper1_wdata_dup_0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y9_2 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p1_int[27]),.T2I1(lint_WDATA_int[27]),.T2I2(nx25587z2),.T2I3(GND),.TB2S(GND),.Q2Z(m0_oper1_wdata_dup_0[27]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y9_3 (.tFragBitInfo(16'b0101010000000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(tcdm_rdata_p1_int[18]),.T3I2(nx25587z2),.T3I3(lint_WDATA_int[18]),.TB3S(GND),.Q3Z(m0_oper1_wdata_dup_0[18]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y10_0 (.tFragBitInfo(16'b0101000101000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(nx25587z2),.T0I2(lint_WDATA_int[21]),.T0I3(tcdm_rdata_p1_int[21]),.TB0S(GND),.Q0Z(m0_oper1_wdata_dup_0[21]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[2]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p1[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y10_2 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[28]),.T2I1(nx25587z2),.T2I2(GND),.T2I3(tcdm_rdata_p1_int[28]),.TB2S(GND),.Q2Z(m0_oper1_wdata_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y10_3 (.tFragBitInfo(16'b0000000010111000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[7]),.T3I1(nx25587z2),.T3I2(tcdm_rdata_p1_int[7]),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper1_wdata_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p1_int[0]),.Q0EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p1[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y11_1 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx36058z2_CAND5_TRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T1I0(m0_oper1_rdata_int[27]),.T1I1(GND),.T1I2(nx11312z1_CAND4_TRSBR_25_tpGCLKBUF),.T1I3(lint_WDATA_int[27]),.TB1S(GND),.Q1Z(tcdm_wdata_p1_dup_0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y11_2 (.tFragBitInfo(16'b0000101000001100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx36058z2_CAND5_TRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[21]),.T2I1(m0_oper1_rdata_int[21]),.T2I2(GND),.T2I3(nx11312z1_CAND4_TRSBR_25_tpGCLKBUF),.TB2S(GND),.Q2Z(tcdm_wdata_p1_dup_0[21]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y11_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y12_0 (.tFragBitInfo(16'b0100110001011111),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T0I0(tcdm_result_p2[22]),.T0I1(tcdm_be_p0_dup_0[2]),.T0I2(NET_106),.T0I3(NET_107),.TB0S(GND),.C0Z(NET_567),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y12_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p1_int[18]),.Q1EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.Q1Z(tcdm_result_p1[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y12_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y12_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y13_0 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_be_p0_17n77s1[2]),.Q0EN(nx40546z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.T0I0(tcdm_addr_p0_dup_0[7]),.T0I1(tcdm_result_p2[7]),.T0I2(NET_107),.T0I3(NET_106),.TB0S(GND),.C0Z(NET_597),.Q0Z(tcdm_be_p1_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y13_1 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx40545z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.T1I0(lint_WDATA_int[22]),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND),.C1Z(tcdm_be_p0_17n77s1[2]),.Q1Z(tcdm_be_p0_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_Y13_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0001001101011111),.B2I0(tcdm_addr_p1_dup_0[7]),.B2I1(NET_114),.B2I2(NET_115),.B2I3(fpgaio_in_int[39]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx40545z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.T2I0(lint_WDATA_int[21]),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND),.B2Z(NET_598),.C2Z(tcdm_be_p0_17n77s1[1]),.Q2Z(tcdm_be_p0_dup_0[1]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_Y13_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_595),.B3I1(NET_596),.B3I2(NET_597),.B3I3(NET_598),.CD3S(VCC),.Q3DI(tcdm_be_p0_17n77s1[1]),.Q3EN(nx40546z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.T3I0(NET_597),.T3I1(NET_598),.T3I2(NET_595),.T3I3(NET_596),.TB3S(NET_599),.C3Z(NET_591),.Q3Z(tcdm_be_p1_dup_0[1]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Y14_0 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000011101110111),.B0I0(NET_114),.B0I1(fpgaio_in_int[38]),.B0I2(tcdm_addr_p1_dup_0[6]),.B0I3(NET_115),.CD0S(GND),.Q0DI(GND),.Q0EN(nx40545z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.T0I0(GND),.T0I1(GND),.T0I2(lint_WDATA_int[20]),.T0I3(GND),.TB0S(GND),.B0Z(NET_798),.C0Z(tcdm_be_p0_17n77s1[0]),.Q0Z(tcdm_be_p0_dup_0[0]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y14_1 (.tFragBitInfo(16'b0001001101011111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_be_p0_17n77s1[3]),.Q1EN(nx40546z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.T1I0(tcdm_addr_p0_dup_0[6]),.T1I1(NET_106),.T1I2(NET_107),.T1I3(tcdm_result_p2[6]),.C1Z(NET_797),.Q1Z(tcdm_be_p1_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Y14_2 (.tFragBitInfo(16'b0000000000000001),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx40545z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(lint_WDATA_int[23]),.TB2S(GND),.C2Z(tcdm_be_p0_17n77s1[3]),.Q2Z(tcdm_be_p0_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_Y14_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_795),.B3I1(NET_797),.B3I2(NET_796),.B3I3(NET_798),.CD3S(VCC),.Q3DI(tcdm_be_p0_17n77s1[0]),.Q3EN(nx40546z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.T3I0(NET_796),.T3I1(NET_798),.T3I2(NET_795),.T3I3(NET_797),.TB3S(NET_799),.C3Z(NET_791),.Q3Z(tcdm_be_p1_dup_0[0]),.B3CO(),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Y15_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y15_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_311),.B1I1(NET_310),.B1I2(NET_312),.B1I3(NET_309),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T1I0(NET_312),.T1I1(NET_309),.T1I2(NET_311),.T1I3(NET_310),.TB1S(NET_313),.C1Z(NET_305),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_Y15_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001001101011111),.B2I0(fpgaio_in_int[44]),.B2I1(NET_115),.B2I2(NET_114),.B2I3(tcdm_addr_p1_dup_0[12]),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[4]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p0_dup_0[12]),.T2I1(NET_107),.T2I2(NET_106),.T2I3(tcdm_result_p2[12]),.TB2S(GND),.B2Z(NET_312),.C2Z(NET_311),.Q2Z(tcdm_result_p1[4]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_Y15_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_be_p0_17n77s1[2]),.Q0EN(nx40547z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_be_p2_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_be_p0_17n77s1[1]),.Q1EN(nx40548z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_be_p3_dup_0[1]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y16_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_be_p0_17n77s1[2]),.Q2EN(nx40548z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_be_p3_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_be_p0_17n77s1[1]),.Q3EN(nx40547z1),.QCK(CLK_int_0__CAND0_TRSBR_25_padClk),.QRT(GND),.QST(GND),.Q3Z(tcdm_be_p2_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y17_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_be_p0_17n77s1[0]),.Q0EN(nx40547z1),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_be_p2_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_be_p0_17n77s1[3]),.Q1EN(nx40548z1),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_be_p3_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_be_p0_17n77s1[3]),.Q2EN(nx40547z1),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(GND),.QST(GND),.Q2Z(tcdm_be_p2_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(GND),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y18_0 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_118),.B0I1(tcdm_addr_p2_dup_0[6]),.B0I2(fpgaio_out_dup_0[70]),.B0I3(NET_104),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.T0I0(nx63842z2_CAND1_BRSTR_25_tpGCLKBUF),.T0I1(GND),.T0I2(GND),.T0I3(RESET_int[0]),.TB0S(GND),.B0Z(NET_796),.C0Z(nx40547z1),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y18_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p2_int[7]),.Q1EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.T1I0(fpgaio_out_dup_0[76]),.T1I1(NET_118),.T1I2(tcdm_addr_p3_dup_0[12]),.T1I3(NET_119),.TB1S(GND),.C1Z(NET_313),.Q1Z(tcdm_result_p2[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_Y18_2 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'b0001010100111111),.B2I0(tcdm_addr_p2_dup_0[12]),.B2I1(i_events[12]),.B2I2(NET_105),.B2I3(NET_104),.CD2S(VCC),.Q2DI(lint_WDATA_int[12]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.T2I0(NET_118),.T2I1(fpgaio_out_dup_0[71]),.T2I2(tcdm_addr_p2_dup_0[7]),.T2I3(NET_104),.TB2S(GND),.B2Z(NET_310),.C2Z(NET_596),.Q2Z(i_events[12]),.B2CO(),.T2CO());

	LOGIC_3 QL_INST_Y18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p2_int[6]),.Q3EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p2[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[31]),.Q0EN(nx40548z1),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(GND),.QST(GND),.Q0Z(tcdm_wen_p3_dup_0),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y19_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_be_p0_17n77s1[0]),.Q1EN(nx40548z1),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(GND),.QST(GND),.Q1Z(tcdm_be_p3_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(GND),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y19_3 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(GND),.QST(GND),.T3I0(nx40548z2_CAND3_BRSTR_25_tpGCLKBUF),.T3I1(GND),.T3I2(RESET_int[0]),.T3I3(GND),.TB3S(GND),.C3Z(nx40548z1),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_Y20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[24]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p3[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y20_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[26]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p3[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y21_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(tcdm_rdata_p2_int[22]),.Q0EN(tcdm_valid_p2_int),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_result_p2[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y21_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y21_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y21_3 (.tFragBitInfo(16'b0000000001111000),.bFragBitInfo(16'b1101111011101110),.B3I0(tcdm_addr_p3_dup_0[10]),.B3I1(nx40548z2_CAND3_BRSTR_25_tpGCLKBUF),.B3I2(NET_201),.B3I3(tcdm_addr_p3_dup_0[9]),.CD3S(GND),.Q3DI(GND),.Q3EN(nx60936z2_CAND5_BRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.T3I0(NET_201),.T3I1(tcdm_addr_p3_dup_0[9]),.T3I2(tcdm_addr_p3_dup_0[10]),.T3I3(nx40548z2_CAND3_BRSTR_25_tpGCLKBUF),.TB3S(lint_WDATA_int[10]),.Q3Z(tcdm_addr_p3_dup_0[10]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y22_0 (.tFragBitInfo(16'b0000000001101100),.bFragBitInfo(16'b1111111101101100),.B0I0(NET_200),.B0I1(tcdm_addr_p3_dup_0[13]),.B0I2(tcdm_addr_p3_dup_0[12]),.B0I3(nx40548z2_CAND3_BRSTR_25_tpGCLKBUF),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60936z2_CAND5_BRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.T0I0(NET_200),.T0I1(tcdm_addr_p3_dup_0[13]),.T0I2(tcdm_addr_p3_dup_0[12]),.T0I3(nx40548z2_CAND3_BRSTR_25_tpGCLKBUF),.TB0S(lint_WDATA_int[13]),.Q0Z(tcdm_addr_p3_dup_0[13]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y22_1 (.tFragBitInfo(16'b0010001000110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx60936z2_CAND5_BRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[14]),.T1I1(GND),.T1I2(NET_199),.T1I3(nx40548z2_CAND3_BRSTR_25_tpGCLKBUF),.TB1S(GND),.Q1Z(tcdm_addr_p3_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y22_2 (.tFragBitInfo(16'b1111000001100110),.bFragBitInfo(16'b1000000000000000),.B2I0(tcdm_addr_p3_dup_0[11]),.B2I1(tcdm_addr_p3_dup_0[10]),.B2I2(NET_201),.B2I3(tcdm_addr_p3_dup_0[9]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx60936z2_CAND5_BRSTR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.T2I0(NET_200),.T2I1(tcdm_addr_p3_dup_0[12]),.T2I2(lint_WDATA_int[12]),.T2I3(nx40548z2_CAND3_BRSTR_25_tpGCLKBUF),.TB2S(GND),.B2Z(NET_200),.Q2Z(tcdm_addr_p3_dup_0[12]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y22_3 (.tFragBitInfo(16'b0111100011110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.T3I0(NET_200),.T3I1(tcdm_addr_p3_dup_0[12]),.T3I2(tcdm_addr_p3_dup_0[14]),.T3I3(tcdm_addr_p3_dup_0[13]),.TB3S(GND),.C3Z(NET_199),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_Y23_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y23_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[20]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[20]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Y23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[3]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p3[3]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y24_0 (.tFragBitInfo(16'b0000101000001100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[10]),.T0I1(tcdm_rdata_p3_int[10]),.T0I2(GND),.T0I3(nx3850z2),.TB0S(GND),.Q0Z(m1_oper1_wdata_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y24_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y24_2 (.tFragBitInfo(16'b0000010100000100),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(NET_0),.T2I2(GND),.T2I3(p3_fsm[2]),.TB2S(GND),.C2Z(nx25788z3),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_Y24_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_25_padClk),.QRT(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y25_0 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx25788z3_CAND4_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[23]),.T0I1(NET_0_CAND1_BRSBR_25_tpGCLKBUF),.T0I2(GND),.T0I3(m1_oper1_rdata_int[23]),.TB0S(GND),.Q0Z(tcdm_wdata_p3_dup_0[23]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y25_1 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx25788z3_CAND4_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T1I0(m1_oper1_rdata_int[29]),.T1I1(GND),.T1I2(NET_0_CAND1_BRSBR_25_tpGCLKBUF),.T1I3(lint_WDATA_int[29]),.TB1S(GND),.Q1Z(tcdm_wdata_p3_dup_0[29]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y25_2 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx3786z2_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_WDATA_int[20]),.T2I2(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.T2I3(tcdm_rdata_p3_int[20]),.TB2S(GND),.Q2Z(m1_oper1_wdata_dup_0[20]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y25_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx3786z2_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[23]),.T3I1(tcdm_rdata_p3_int[23]),.T3I2(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper1_wdata_dup_0[23]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y26_0 (.tFragBitInfo(16'b0101010000000100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx25788z3_CAND4_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(m1_oper1_rdata_int[30]),.T0I2(NET_0_CAND1_BRSBR_25_tpGCLKBUF),.T0I3(lint_WDATA_int[30]),.TB0S(GND),.Q0Z(tcdm_wdata_p3_dup_0[30]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y26_1 (.tFragBitInfo(16'b0100010001010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx25788z3_CAND4_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(lint_WDATA_int[31]),.T1I2(m1_oper1_rdata_int[31]),.T1I3(NET_0_CAND1_BRSBR_25_tpGCLKBUF),.TB1S(GND),.Q1Z(tcdm_wdata_p3_dup_0[31]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y26_2 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx3786z2_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.T2I1(lint_WDATA_int[18]),.T2I2(GND),.T2I3(tcdm_rdata_p3_int[18]),.TB2S(GND),.Q2Z(m1_oper1_wdata_dup_0[18]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y26_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx25788z3_CAND4_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[21]),.T3I1(m1_oper1_rdata_int[21]),.T3I2(NET_0_CAND1_BRSBR_25_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p3_dup_0[21]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y27_0 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx25788z3_CAND4_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T0I0(NET_0_CAND1_BRSBR_25_tpGCLKBUF),.T0I1(GND),.T0I2(lint_WDATA_int[27]),.T0I3(m1_oper1_rdata_int[27]),.TB0S(GND),.Q0Z(tcdm_wdata_p3_dup_0[27]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y27_1 (.tFragBitInfo(16'b0000110000001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx3786z2_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p3_int[27]),.T1I1(lint_WDATA_int[27]),.T1I2(GND),.T1I3(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.TB1S(GND),.Q1Z(m1_oper1_wdata_dup_0[27]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y27_2 (.tFragBitInfo(16'b0011001000010000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx25788z3_CAND4_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(NET_0_CAND1_BRSBR_25_tpGCLKBUF),.T2I1(GND),.T2I2(m1_oper1_rdata_int[28]),.T2I3(lint_WDATA_int[28]),.TB2S(GND),.Q2Z(tcdm_wdata_p3_dup_0[28]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y27_3 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx3786z2_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T3I0(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.T3I1(tcdm_rdata_p3_int[24]),.T3I2(lint_WDATA_int[24]),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper1_wdata_dup_0[24]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y28_0 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx3786z2_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[22]),.T0I1(GND),.T0I2(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.T0I3(tcdm_rdata_p3_int[22]),.TB0S(GND),.Q0Z(m1_oper1_wdata_dup_0[22]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y28_1 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx3786z2_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T1I0(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.T1I1(lint_WDATA_int[28]),.T1I2(tcdm_rdata_p3_int[28]),.T1I3(GND),.TB1S(GND),.Q1Z(m1_oper1_wdata_dup_0[28]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y28_2 (.tFragBitInfo(16'b0000111000000100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx3786z2_CAND5_BRSBR_25_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.T2I1(tcdm_rdata_p3_int[26]),.T2I2(GND),.T2I3(lint_WDATA_int[26]),.TB2S(GND),.Q2Z(m1_oper1_wdata_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y28_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y29_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T0I0(NET_303),.T0I1(m1_oper1_waddr_dup_0[6]),.T0I2(m1_oper1_waddr_dup_0[7]),.T0I3(m1_oper1_waddr_dup_0[8]),.TB0S(GND),.C0Z(NET_671),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y29_1 (.tFragBitInfo(16'b1010000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[8]),.T1I1(NET_744),.T1I2(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.T1I3(p3_fsm[0]),.TB1S(GND),.Q1Z(m1_oper1_waddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y29_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0111111110000000),.B2I0(NET_303),.B2I1(m1_oper1_waddr_dup_0[6]),.B2I2(m1_oper1_waddr_dup_0[7]),.B2I3(m1_oper1_waddr_dup_0[8]),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_waddr_dup_0[5]),.T2I1(m1_oper1_waddr_dup_0[3]),.T2I2(m1_oper1_waddr_dup_0[4]),.T2I3(m1_oper1_waddr_dup_0[2]),.TB2S(GND),.B2Z(NET_744),.C2Z(NET_303),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_Y29_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Y30_0 (.tFragBitInfo(16'b0111100011110000),.bFragBitInfo(16'b0000010000000001),.B0I0(m1_oper1_waddr_dup_0[10]),.B0I1(m1_oper1_waddr_dup_0[8]),.B0I2(m1_oper1_waddr_dup_0[11]),.B0I3(control_in_int[22]),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_waddr_dup_0[10]),.T0I1(NET_671),.T0I2(m1_oper1_waddr_dup_0[11]),.T0I3(m1_oper1_waddr_dup_0[9]),.TB0S(GND),.B0Z(NET_226),.C0Z(NET_692),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y30_1 (.tFragBitInfo(16'b1111000001000100),.bFragBitInfo(16'b1000100010001011),.B1I0(lint_ADDR_int[9]),.B1I1(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.B1I2(p3_fsm[0]),.B1I3(NET_671),.CD1S(GND),.Q1DI(GND),.Q1EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T1I0(p3_fsm[0]),.T1I1(NET_671),.T1I2(lint_ADDR_int[9]),.T1I3(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.TB1S(m1_oper1_waddr_dup_0[9]),.Q1Z(m1_oper1_waddr_dup_0[9]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y30_2 (.tFragBitInfo(16'b1100110000000101),.bFragBitInfo(16'b0000100100000101),.B2I0(m1_oper1_waddr_dup_0[10]),.B2I1(NET_671),.B2I2(GND),.B2I3(m1_oper1_waddr_dup_0[9]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(p3_fsm[0]),.T2I1(lint_ADDR_int[10]),.T2I2(NET_670),.T2I3(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.TB2S(GND),.B2Z(NET_670),.Q2Z(m1_oper1_waddr_dup_0[10]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y30_3 (.tFragBitInfo(16'b1111000001000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx64401z2),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T3I0(p3_fsm[0]),.T3I1(NET_692),.T3I2(lint_ADDR_int[11]),.T3I3(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF),.TB3S(GND),.Q3Z(m1_oper1_waddr_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y31_0 (.tFragBitInfo(16'b1100101011000000),.bFragBitInfo(16'b0110101010101010),.B0I0(m1_oper1_raddr_dup_0[11]),.B0I1(m1_oper1_raddr_dup_0[10]),.B0I2(m1_oper1_raddr_dup_0[9]),.B0I3(NET_652),.CD0S(GND),.Q0DI(GND),.Q0EN(nx36808z2),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T0I0(p3_fsm[2]),.T0I1(lint_ADDR_int[11]),.T0I2(NET_508),.T0I3(NET_822),.TB0S(GND),.B0Z(NET_822),.Q0Z(m1_oper1_raddr_dup_0[11]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Y31_1 (.tFragBitInfo(16'b1100101011000000),.bFragBitInfo(16'b1011101000010000),.B1I0(NET_508),.B1I1(NET_652),.B1I2(p3_fsm[2]),.B1I3(lint_ADDR_int[9]),.CD1S(GND),.Q1DI(GND),.Q1EN(nx36808z2),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T1I0(p3_fsm[2]),.T1I1(lint_ADDR_int[9]),.T1I2(NET_508),.T1I3(NET_652),.TB1S(m1_oper1_raddr_dup_0[9]),.Q1Z(m1_oper1_raddr_dup_0[9]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Y31_2 (.tFragBitInfo(16'b1010111000000100),.bFragBitInfo(16'b0010000100010001),.B2I0(m1_oper1_raddr_dup_0[10]),.B2I1(GND),.B2I2(m1_oper1_raddr_dup_0[9]),.B2I3(NET_652),.CD2S(GND),.Q2DI(GND),.Q2EN(nx36808z2),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T2I0(NET_508),.T2I1(p3_fsm[2]),.T2I2(NET_821),.T2I3(lint_ADDR_int[10]),.TB2S(GND),.B2Z(NET_821),.Q2Z(m1_oper1_raddr_dup_0[10]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Y31_3 (.tFragBitInfo(16'b1110010010100000),.bFragBitInfo(16'b1010000010101100),.B3I0(lint_ADDR_int[3]),.B3I1(p3_fsm[2]),.B3I2(NET_508),.B3I3(m1_oper1_raddr_dup_0[2]),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36808z2),.QCK(CLK_int_0__CAND0_BRSBR_25_padClk),.QRT(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF),.QST(GND),.T3I0(NET_508),.T3I1(m1_oper1_raddr_dup_0[2]),.T3I2(lint_ADDR_int[3]),.T3I3(p3_fsm[2]),.TB3S(m1_oper1_raddr_dup_0[3]),.Q3Z(m1_oper1_raddr_dup_0[3]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Y32_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Y32_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Y32_2 (.tFragBitInfo(16'b0000011000001010),.bFragBitInfo(16'b0000000000000000),.T2I0(m1_oper1_raddr_dup_0[4]),.T2I1(m1_oper1_raddr_dup_0[3]),.T2I2(GND),.T2I3(m1_oper1_raddr_dup_0[2]),.TB2S(GND),.C2Z(NET_530),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_Y32_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z1_0 (.tFragBitInfo(16'b0000000000001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T0I1(lint_ADDR_int[1]),.T0I2(GND),.T0I3(GND),.TB0S(GND),.Q0Z(m0_oper1_waddr_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z1_1 (.tFragBitInfo(16'b0000001000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[0]),.T1I1(GND),.T1I2(GND),.T1I3(NET_77),.TB1S(GND),.Q1Z(m0_oper1_raddr_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z1_2 (.tFragBitInfo(16'b0000000000100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[0]),.T2I1(GND),.T2I2(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T2I3(GND),.TB2S(GND),.Q2Z(m0_oper1_waddr_dup_0[0]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z1_3 (.tFragBitInfo(16'b0000010000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(lint_ADDR_int[1]),.T3I2(GND),.T3I3(NET_77),.TB3S(GND),.Q3Z(m0_oper1_raddr_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z2_0 (.tFragBitInfo(16'b1100101011000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(p1_cnt[6]),.T0I1(lint_ADDR_int[8]),.T0I2(NET_77),.T0I3(p1_fsm[4]),.TB0S(GND),.Q0Z(m0_oper1_raddr_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z2_1 (.tFragBitInfo(16'b1100101011000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(p1_cnt[4]),.T1I1(lint_ADDR_int[6]),.T1I2(NET_77),.T1I3(p1_fsm[4]),.TB1S(GND),.Q1Z(m0_oper1_raddr_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z2_2 (.tFragBitInfo(16'b1100110010100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(p1_cnt[6]),.T2I1(lint_ADDR_int[8]),.T2I2(p1_fsm[3]),.T2I3(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.TB2S(GND),.Q2Z(m0_oper1_waddr_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z2_3 (.tFragBitInfo(16'b1100110010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(p1_cnt[4]),.T3I1(lint_ADDR_int[6]),.T3I2(p1_fsm[3]),.T3I3(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.TB3S(GND),.Q3Z(m0_oper1_waddr_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z3_0 (.tFragBitInfo(16'b1110001011000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(p1_cnt[3]),.T0I1(NET_77),.T0I2(lint_ADDR_int[5]),.T0I3(p1_fsm[4]),.TB0S(GND),.Q0Z(m0_oper1_raddr_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z3_1 (.tFragBitInfo(16'b1111100000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(p1_cnt[0]),.T1I1(p1_fsm[3]),.T1I2(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T1I3(lint_ADDR_int[2]),.TB1S(GND),.Q1Z(m0_oper1_waddr_dup_0[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z3_2 (.tFragBitInfo(16'b1110010010100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx18281z3),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(NET_77),.T2I1(p1_cnt[0]),.T2I2(lint_ADDR_int[2]),.T2I3(p1_fsm[4]),.TB2S(GND),.Q2Z(m0_oper1_raddr_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z3_3 (.tFragBitInfo(16'b1111100000001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx35588z2),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(p1_cnt[3]),.T3I1(p1_fsm[3]),.T3I2(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T3I3(lint_ADDR_int[5]),.TB3S(GND),.Q3Z(m0_oper1_waddr_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z4_0 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx36058z2_CAND4_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[24]),.T0I1(nx11312z1_CAND3_TRSTR_26_tpGCLKBUF),.T0I2(GND),.T0I3(m0_oper1_rdata_int[24]),.TB0S(GND),.Q0Z(tcdm_wdata_p1_dup_0[24]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z4_1 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx36058z2_CAND4_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[19]),.T1I1(m0_oper1_rdata_int[19]),.T1I2(nx11312z1_CAND3_TRSTR_26_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p1_dup_0[19]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z4_2 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx36058z2_CAND4_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(nx11312z1_CAND3_TRSTR_26_tpGCLKBUF),.T2I1(GND),.T2I2(lint_WDATA_int[26]),.T2I3(m0_oper1_rdata_int[26]),.TB2S(GND),.Q2Z(tcdm_wdata_p1_dup_0[26]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z4_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z5_0 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[10]),.T0I1(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T0I2(GND),.T0I3(tcdm_rdata_p1_int[10]),.TB0S(GND),.Q0Z(m0_oper1_wdata_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z5_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p1_int[11]),.T1I1(lint_WDATA_int[11]),.T1I2(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(m0_oper1_wdata_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z5_2 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T2I1(GND),.T2I2(lint_WDATA_int[8]),.T2I3(tcdm_rdata_p1_int[8]),.TB2S(GND),.Q2Z(m0_oper1_wdata_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z5_3 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p1_int[5]),.T3I1(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T3I2(lint_WDATA_int[5]),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper1_wdata_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z6_1 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p1_int[3]),.T1I1(GND),.T1I2(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T1I3(lint_WDATA_int[3]),.TB1S(GND),.Q1Z(m0_oper1_wdata_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z6_2 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p1_int[2]),.T2I1(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T2I2(lint_WDATA_int[2]),.T2I3(GND),.TB2S(GND),.Q2Z(m0_oper1_wdata_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z6_3 (.tFragBitInfo(16'b0101000101000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T3I2(lint_WDATA_int[9]),.T3I3(tcdm_rdata_p1_int[9]),.TB3S(GND),.Q3Z(m0_oper1_wdata_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_716),.B0I1(tcdm_addr_p0_dup_0[6]),.B0I2(tcdm_addr_p0_dup_0[8]),.B0I3(tcdm_addr_p0_dup_0[7]),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.B0Z(NET_737),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z7_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p0_dup_0[9]),.T1I1(tcdm_addr_p0_dup_0[10]),.T1I2(tcdm_addr_p0_dup_0[11]),.T1I3(NET_737),.C1Z(NET_788),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Z7_2 (.tFragBitInfo(16'b1100010111001010),.bFragBitInfo(16'b0111100011110000),.B2I0(tcdm_addr_p0_dup_0[9]),.B2I1(tcdm_addr_p0_dup_0[10]),.B2I2(tcdm_addr_p0_dup_0[11]),.B2I3(NET_737),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p0_dup_0[9]),.T2I1(lint_WDATA_int[9]),.T2I2(nx45272z2),.T2I3(NET_737),.TB2S(GND),.B2Z(NET_815),.Q2Z(tcdm_addr_p0_dup_0[9]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z7_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[11]),.T3I1(NET_815),.T3I2(nx45272z2),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_addr_p0_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z8_0 (.tFragBitInfo(16'b0000111000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p1_int[0]),.T0I1(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T0I2(GND),.T0I3(lint_WDATA_int[0]),.TB0S(GND),.Q0Z(m0_oper1_wdata_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z8_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(tcdm_rdata_p1_int[17]),.T1I1(lint_WDATA_int[17]),.T1I2(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(m0_oper1_wdata_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z8_2 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[12]),.T2I1(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T2I2(GND),.T2I3(tcdm_rdata_p1_int[12]),.TB2S(GND),.Q2Z(m0_oper1_wdata_dup_0[12]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z8_3 (.tFragBitInfo(16'b0000000010111000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_26_padClk),.QRT(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[1]),.T3I1(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF),.T3I2(tcdm_rdata_p1_int[1]),.T3I3(GND),.TB3S(GND),.Q3Z(m0_oper1_wdata_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z9_0 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p1_int[13]),.T0I1(nx25587z2),.T0I2(lint_WDATA_int[13]),.T0I3(GND),.TB0S(GND),.Q0Z(m0_oper1_wdata_dup_0[13]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z9_1 (.tFragBitInfo(16'b0011001100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(tcdm_req_p1_dup_0),.T1I1(GND),.T1I2(p1_fsm[4]),.T1I3(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF),.TB1S(GND),.C1Z(nx13970z2),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_Z9_2 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p1_int[14]),.T2I1(nx25587z2),.T2I2(lint_WDATA_int[14]),.T2I3(GND),.TB2S(GND),.Q2Z(m0_oper1_wdata_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z9_3 (.tFragBitInfo(16'b0101010000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(nx25587z2),.T3I2(tcdm_rdata_p1_int[4]),.T3I3(lint_WDATA_int[4]),.TB3S(GND),.Q3Z(m0_oper1_wdata_dup_0[4]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z10_0 (.tFragBitInfo(16'b0000101000001100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[15]),.T0I1(tcdm_rdata_p1_int[15]),.T0I2(GND),.T0I3(nx25587z2),.TB0S(GND),.Q0Z(m0_oper1_wdata_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z10_1 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx36058z2_CAND5_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[25]),.T1I1(GND),.T1I2(nx11312z1_CAND4_TRSBR_26_tpGCLKBUF),.T1I3(m0_oper1_rdata_int[25]),.TB1S(GND),.Q1Z(tcdm_wdata_p1_dup_0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z10_2 (.tFragBitInfo(16'b0101000001000100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(tcdm_rdata_p1_int[16]),.T2I2(lint_WDATA_int[16]),.T2I3(nx25587z2),.TB2S(GND),.Q2Z(m0_oper1_wdata_dup_0[16]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z10_3 (.tFragBitInfo(16'b0000110000001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx39177z2),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p1_int[6]),.T3I1(lint_WDATA_int[6]),.T3I2(GND),.T3I3(nx25587z2),.TB3S(GND),.Q3Z(m0_oper1_wdata_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z11_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[1]),.Q0EN(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p1_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z11_1 (.tFragBitInfo(16'b0011001000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx36058z2_CAND5_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(nx11312z1_CAND4_TRSBR_26_tpGCLKBUF),.T1I1(GND),.T1I2(m0_oper1_rdata_int[20]),.T1I3(lint_WDATA_int[20]),.TB1S(GND),.Q1Z(tcdm_wdata_p1_dup_0[20]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z11_2 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx36058z2_CAND5_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T2I0(nx11312z1_CAND4_TRSBR_26_tpGCLKBUF),.T2I1(lint_WDATA_int[22]),.T2I2(GND),.T2I3(m0_oper1_rdata_int[22]),.TB2S(GND),.Q2Z(tcdm_wdata_p1_dup_0[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z11_3 (.tFragBitInfo(16'b0000000010001011),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx13970z2_CAND2_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[2]),.T3I1(NET_89),.T3I2(tcdm_addr_p1_dup_0[2]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_addr_p1_dup_0[2]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z12_0 (.tFragBitInfo(16'b0000000001101010),.bFragBitInfo(16'b1101111011101110),.B0I0(tcdm_addr_p1_dup_0[17]),.B0I1(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF),.B0I2(tcdm_addr_p1_dup_0[16]),.B0I3(NET_327),.CD0S(GND),.Q0DI(GND),.Q0EN(nx13970z2_CAND2_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T0I0(tcdm_addr_p1_dup_0[17]),.T0I1(NET_327),.T0I2(tcdm_addr_p1_dup_0[16]),.T0I3(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF),.TB0S(lint_WDATA_int[17]),.Q0Z(tcdm_addr_p1_dup_0[17]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z12_1 (.tFragBitInfo(16'b1010101000111100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx13970z2_CAND2_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[16]),.T1I1(NET_327),.T1I2(tcdm_addr_p1_dup_0[16]),.T1I3(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF),.TB1S(GND),.Q1Z(tcdm_addr_p1_dup_0[16]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z12_2 (.tFragBitInfo(16'b1100110001011010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx13970z2_CAND2_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p1_dup_0[19]),.T2I1(lint_WDATA_int[19]),.T2I2(NET_326),.T2I3(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF),.TB2S(GND),.Q2Z(tcdm_addr_p1_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z12_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p1_int[16]),.Q3EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(tcdm_addr_p1_dup_0[18]),.T3I1(tcdm_addr_p1_dup_0[17]),.T3I2(tcdm_addr_p1_dup_0[16]),.T3I3(NET_327),.TB3S(GND),.C3Z(NET_326),.Q3Z(tcdm_result_p1[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_Z13_0 (.tFragBitInfo(16'b1011000111100100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx13970z2_CAND2_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T0I0(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF),.T0I1(NET_350),.T0I2(lint_WDATA_int[18]),.T0I3(tcdm_addr_p1_dup_0[18]),.TB0S(GND),.Q0Z(tcdm_addr_p1_dup_0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z13_1 (.tFragBitInfo(16'b1011111000010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx13970z2_CAND2_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF),.T1I1(NET_351),.T1I2(tcdm_addr_p1_dup_0[12]),.T1I3(lint_WDATA_int[12]),.TB1S(GND),.Q1Z(tcdm_addr_p1_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z13_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_352),.B2I1(tcdm_addr_p1_dup_0[16]),.B2I2(NET_351),.B2I3(tcdm_addr_p1_dup_0[15]),.CD2S(VCC),.Q2DI(tcdm_rdata_p1_int[14]),.Q2EN(tcdm_valid_p1_int),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T2I0(NET_352),.T2I1(tcdm_addr_p1_dup_0[16]),.T2I2(NET_351),.T2I3(tcdm_addr_p1_dup_0[15]),.TB2S(tcdm_addr_p1_dup_0[17]),.C2Z(NET_350),.Q2Z(tcdm_result_p1[14]),.B2CO(),.B2Z(),.T2CO());

	LOGIC_3 QL_INST_Z13_3 (.tFragBitInfo(16'b0000011100001000),.bFragBitInfo(16'b1011111011101110),.B3I0(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF),.B3I1(tcdm_addr_p1_dup_0[15]),.B3I2(NET_352),.B3I3(NET_351),.CD3S(GND),.Q3DI(GND),.Q3EN(nx13970z2_CAND2_TRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(NET_352),.T3I1(NET_351),.T3I2(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF),.T3I3(tcdm_addr_p1_dup_0[15]),.TB3S(lint_WDATA_int[15]),.Q3Z(tcdm_addr_p1_dup_0[15]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z14_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z14_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[13]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(NET_50),.T1I1(tcdm_addr_p1_dup_0[13]),.T1I2(i_events[13]),.T1I3(NET_51),.C1Z(NET_347),.Q1Z(i_events[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Z14_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(lint_WDATA_int[5]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.Q2Z(i_events[5]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z14_3 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_26_padClk),.QRT(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(NET_50),.T3I1(tcdm_addr_p1_dup_0[5]),.T3I2(i_events[5]),.T3I3(NET_51),.C3Z(NET_835),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_Z17_0 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx63842z2_CAND1_BRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(tcdm_addr_p2_dup_0[11]),.T0I1(NET_51),.T0I2(i_events[11]),.T0I3(NET_253),.TB0S(GND),.C0Z(NET_299),.Q0Z(tcdm_addr_p2_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z17_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[2]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.Q1Z(i_events[2]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z17_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001010100111111),.B2I0(NET_105),.B2I1(tcdm_addr_p2_dup_0[2]),.B2I2(NET_104),.B2I3(i_events[2]),.CD2S(VCC),.Q2DI(lint_WDATA_int[11]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.B2Z(NET_898),.Q2Z(i_events[11]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z17_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z18_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[7]),.Q1EN(nx60509z1),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(NET_119),.T1I1(tcdm_addr_p3_dup_0[7]),.T1I2(i_events[7]),.T1I3(NET_105),.TB1S(GND),.C1Z(NET_599),.Q1Z(i_events[7]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_Z18_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_119),.B2I1(i_events[6]),.B2I2(tcdm_addr_p3_dup_0[6]),.B2I3(NET_105),.CD2S(VCC),.Q2DI(lint_WDATA_int[6]),.Q2EN(nx60509z1),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.B2Z(NET_799),.Q2Z(i_events[6]),.B2CO(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z18_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0001001101011111),.B0I0(NET_104),.B0I1(NET_119),.B0I2(tcdm_addr_p2_dup_0[17]),.B0I3(tcdm_addr_p3_dup_0[17]),.B0Z(NET_445),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z19_1 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.T1I0(NET_104),.T1I1(tcdm_addr_p3_dup_0[19]),.T1I2(NET_119),.T1I3(tcdm_addr_p2_dup_0[19]),.C1Z(NET_493),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Z19_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_Z20_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z20_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z20_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD2S(VCC),.Q2DI(tcdm_rdata_p3_int[2]),.Q2EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.Q2Z(tcdm_result_p3[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z20_3 (.tFragBitInfo(16'b0000000000110101),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(tcdm_addr_p2_dup_0[18]),.T3I1(tcdm_addr_p3_dup_0[18]),.T3I2(lint_ADDR_int[2]),.T3I3(GND),.TB3S(GND),.C3Z(NET_472),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_Z21_0 (.tFragBitInfo(16'b0000111000000100),.bFragBitInfo(16'b1000000000000000),.B0I0(tcdm_addr_p3_dup_0[17]),.B0I1(tcdm_addr_p3_dup_0[16]),.B0I2(tcdm_addr_p3_dup_0[15]),.B0I3(NET_301),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60936z2_CAND5_BRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(nx40548z2_CAND3_BRSTR_26_tpGCLKBUF),.T0I1(NET_847),.T0I2(GND),.T0I3(lint_WDATA_int[17]),.TB0S(GND),.B0Z(NET_846),.Q0Z(tcdm_addr_p3_dup_0[17]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z21_1 (.tFragBitInfo(16'b1011111000010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx60936z2_CAND5_BRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(nx40548z2_CAND3_BRSTR_26_tpGCLKBUF),.T1I1(NET_846),.T1I2(tcdm_addr_p3_dup_0[18]),.T1I3(lint_WDATA_int[18]),.TB1S(GND),.Q1Z(tcdm_addr_p3_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z21_2 (.tFragBitInfo(16'b0000100000000000),.bFragBitInfo(16'b0110101010101010),.B2I0(tcdm_addr_p3_dup_0[17]),.B2I1(tcdm_addr_p3_dup_0[16]),.B2I2(tcdm_addr_p3_dup_0[15]),.B2I3(NET_301),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p3_dup_0[13]),.T2I1(tcdm_addr_p3_dup_0[14]),.T2I2(GND),.T2I3(tcdm_addr_p3_dup_0[12]),.TB2S(GND),.B2Z(NET_847),.C2Z(NET_302),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_Z21_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(NET_201),.B3I1(tcdm_addr_p3_dup_0[10]),.B3I2(tcdm_addr_p3_dup_0[11]),.B3I3(NET_302),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(tcdm_addr_p3_dup_0[11]),.T3I1(NET_302),.T3I2(NET_201),.T3I3(tcdm_addr_p3_dup_0[10]),.TB3S(tcdm_addr_p3_dup_0[9]),.C3Z(NET_301),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_Z22_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0110101010101010),.B0I0(tcdm_addr_p3_dup_0[11]),.B0I1(NET_201),.B0I2(tcdm_addr_p3_dup_0[9]),.B0I3(tcdm_addr_p3_dup_0[10]),.CD0S(VCC),.Q0DI(tcdm_rdata_p3_int[13]),.Q0EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(tcdm_addr_p3_dup_0[8]),.T0I1(NET_202),.T0I2(tcdm_addr_p3_dup_0[6]),.T0I3(tcdm_addr_p3_dup_0[7]),.TB0S(GND),.B0Z(NET_631),.C0Z(NET_201),.Q0Z(tcdm_result_p3[13]),.B0CO(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z22_1 (.tFragBitInfo(16'b1011111000010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx60936z2_CAND5_BRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(nx40548z2_CAND3_BRSTR_26_tpGCLKBUF),.T1I1(NET_201),.T1I2(tcdm_addr_p3_dup_0[9]),.T1I3(lint_WDATA_int[9]),.TB1S(GND),.Q1Z(tcdm_addr_p3_dup_0[9]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z22_2 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx60936z2_CAND5_BRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(nx40548z2_CAND3_BRSTR_26_tpGCLKBUF),.T2I1(lint_WDATA_int[11]),.T2I2(GND),.T2I3(NET_631),.TB2S(GND),.Q2Z(tcdm_addr_p3_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z22_3 (.tFragBitInfo(16'b1000110111011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx60936z2_CAND5_BRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(nx40548z2_CAND3_BRSTR_26_tpGCLKBUF),.T3I1(lint_WDATA_int[6]),.T3I2(tcdm_addr_p3_dup_0[6]),.T3I3(NET_202),.TB3S(GND),.Q3Z(tcdm_addr_p3_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z23_0 (.tFragBitInfo(16'b0000000001101010),.bFragBitInfo(16'b1111111101101010),.B0I0(tcdm_addr_p3_dup_0[7]),.B0I1(tcdm_addr_p3_dup_0[6]),.B0I2(NET_202),.B0I3(nx40548z2_CAND3_BRSTR_26_tpGCLKBUF),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60936z2_CAND5_BRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(tcdm_addr_p3_dup_0[7]),.T0I1(tcdm_addr_p3_dup_0[6]),.T0I2(NET_202),.T0I3(nx40548z2_CAND3_BRSTR_26_tpGCLKBUF),.TB0S(lint_WDATA_int[7]),.Q0Z(tcdm_addr_p3_dup_0[7]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z23_1 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(tcdm_rdata_p3_int[8]),.Q1EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p3_dup_0[3]),.T1I1(tcdm_addr_p3_dup_0[2]),.T1I2(tcdm_addr_p3_dup_0[4]),.T1I3(tcdm_addr_p3_dup_0[5]),.TB1S(GND),.C1Z(NET_202),.Q1Z(tcdm_result_p3[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_Z23_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0111111110000000),.B2I0(tcdm_addr_p3_dup_0[7]),.B2I1(tcdm_addr_p3_dup_0[6]),.B2I2(NET_202),.B2I3(tcdm_addr_p3_dup_0[8]),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.B2Z(NET_816),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z23_3 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx60936z2_CAND5_BRSTR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(NET_816),.T3I1(nx40548z2_CAND3_BRSTR_26_tpGCLKBUF),.T3I2(lint_WDATA_int[8]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_addr_p3_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z24_0 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T0I0(nx3850z2),.T0I1(lint_WDATA_int[1]),.T0I2(GND),.T0I3(tcdm_rdata_p3_int[1]),.TB0S(GND),.Q0Z(m1_oper1_wdata_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z24_1 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T1I0(nx3850z2),.T1I1(tcdm_rdata_p3_int[11]),.T1I2(lint_WDATA_int[11]),.T1I3(GND),.TB1S(GND),.Q1Z(m1_oper1_wdata_dup_0[11]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z24_2 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T2I0(tcdm_rdata_p3_int[4]),.T2I1(GND),.T2I2(nx3850z2),.T2I3(lint_WDATA_int[4]),.TB2S(GND),.Q2Z(m1_oper1_wdata_dup_0[4]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z24_3 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSTR_26_padClk),.QRT(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF),.QST(GND),.T3I0(nx3850z2),.T3I1(tcdm_rdata_p3_int[9]),.T3I2(lint_WDATA_int[9]),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper1_wdata_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z25_0 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx3786z2_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T0I0(nx3850z2_CAND3_BRSBR_26_tpGCLKBUF),.T0I1(lint_WDATA_int[8]),.T0I2(GND),.T0I3(tcdm_rdata_p3_int[8]),.TB0S(GND),.Q0Z(m1_oper1_wdata_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z25_1 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx3786z2_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(nx3850z2_CAND3_BRSBR_26_tpGCLKBUF),.T1I1(lint_WDATA_int[0]),.T1I2(GND),.T1I3(tcdm_rdata_p3_int[0]),.TB1S(GND),.Q1Z(m1_oper1_wdata_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z25_2 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx3786z2_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T2I0(nx3850z2_CAND3_BRSBR_26_tpGCLKBUF),.T2I1(lint_WDATA_int[14]),.T2I2(GND),.T2I3(tcdm_rdata_p3_int[14]),.TB2S(GND),.Q2Z(m1_oper1_wdata_dup_0[14]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z25_3 (.tFragBitInfo(16'b0010001000110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx3786z2_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[13]),.T3I1(GND),.T3I2(tcdm_rdata_p3_int[13]),.T3I3(nx3850z2_CAND3_BRSBR_26_tpGCLKBUF),.TB3S(GND),.Q3Z(m1_oper1_wdata_dup_0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z26_0 (.tFragBitInfo(16'b0000110000001010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx3786z2_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T0I0(tcdm_rdata_p3_int[17]),.T0I1(lint_WDATA_int[17]),.T0I2(GND),.T0I3(nx3850z2_CAND3_BRSBR_26_tpGCLKBUF),.TB0S(GND),.Q0Z(m1_oper1_wdata_dup_0[17]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z26_1 (.tFragBitInfo(16'b0010001000110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx3786z2_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[6]),.T1I1(GND),.T1I2(tcdm_rdata_p3_int[6]),.T1I3(nx3850z2_CAND3_BRSBR_26_tpGCLKBUF),.TB1S(GND),.Q1Z(m1_oper1_wdata_dup_0[6]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z26_2 (.tFragBitInfo(16'b0000101100001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx25788z3_CAND4_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[22]),.T2I1(NET_0_CAND1_BRSBR_26_tpGCLKBUF),.T2I2(GND),.T2I3(m1_oper1_rdata_int[22]),.TB2S(GND),.Q2Z(tcdm_wdata_p3_dup_0[22]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z26_3 (.tFragBitInfo(16'b0000000010111000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx25788z3_CAND4_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[20]),.T3I1(NET_0_CAND1_BRSBR_26_tpGCLKBUF),.T3I2(m1_oper1_rdata_int[20]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p3_dup_0[20]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z27_0 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx3786z2_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(lint_WDATA_int[12]),.T0I2(nx3850z2_CAND3_BRSBR_26_tpGCLKBUF),.T0I3(tcdm_rdata_p3_int[12]),.TB0S(GND),.Q0Z(m1_oper1_wdata_dup_0[12]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z27_1 (.tFragBitInfo(16'b0000110000001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx25788z3_CAND4_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(m1_oper1_rdata_int[25]),.T1I1(lint_WDATA_int[25]),.T1I2(GND),.T1I3(NET_0_CAND1_BRSBR_26_tpGCLKBUF),.TB1S(GND),.Q1Z(tcdm_wdata_p3_dup_0[25]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z27_2 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx25788z3_CAND4_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_rdata_int[24]),.T2I1(lint_WDATA_int[24]),.T2I2(NET_0_CAND1_BRSBR_26_tpGCLKBUF),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_wdata_p3_dup_0[24]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z27_3 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx25788z3_CAND4_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(m1_oper1_rdata_int[26]),.T3I1(NET_0_CAND1_BRSBR_26_tpGCLKBUF),.T3I2(lint_WDATA_int[26]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p3_dup_0[26]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z28_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_Z28_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_Z28_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_Z28_3 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx3786z2_CAND5_BRSBR_26_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(tcdm_rdata_p3_int[16]),.T3I1(nx3850z2_CAND3_BRSBR_26_tpGCLKBUF),.T3I2(lint_WDATA_int[16]),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper1_wdata_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z30_0 (.tFragBitInfo(16'b1101110000010000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx36808z2),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_raddr_dup_0[2]),.T0I1(NET_508),.T0I2(p3_fsm[2]),.T0I3(lint_ADDR_int[2]),.TB0S(GND),.Q0Z(m1_oper1_raddr_dup_0[2]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z30_1 (.tFragBitInfo(16'b0000000001101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(NET_572),.T1I1(m1_oper1_raddr_dup_0[7]),.T1I2(m1_oper1_raddr_dup_0[6]),.T1I3(GND),.C1Z(NET_613),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_Z30_2 (.tFragBitInfo(16'b1011100010001000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx36808z2),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T2I0(lint_ADDR_int[7]),.T2I1(NET_508),.T2I2(NET_613),.T2I3(p3_fsm[2]),.TB2S(GND),.Q2Z(m1_oper1_raddr_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_Z30_3 (.tFragBitInfo(16'b1110001011000000),.bFragBitInfo(16'b1010101000001100),.B3I0(lint_ADDR_int[6]),.B3I1(p3_fsm[2]),.B3I2(NET_572),.B3I3(NET_508),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36808z2),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(NET_572),.T3I1(NET_508),.T3I2(lint_ADDR_int[6]),.T3I3(p3_fsm[2]),.TB3S(m1_oper1_raddr_dup_0[6]),.Q3Z(m1_oper1_raddr_dup_0[6]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_Z31_0 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0111100011110000),.B0I0(m1_oper1_raddr_dup_0[7]),.B0I1(m1_oper1_raddr_dup_0[6]),.B0I2(m1_oper1_raddr_dup_0[8]),.B0I3(NET_572),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_raddr_dup_0[3]),.T0I1(m1_oper1_raddr_dup_0[2]),.T0I2(m1_oper1_raddr_dup_0[4]),.T0I3(m1_oper1_raddr_dup_0[5]),.TB0S(GND),.B0Z(NET_632),.C0Z(NET_572),.B0CO(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_Z31_1 (.tFragBitInfo(16'b1010110010100000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx36808z2),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T1I0(lint_ADDR_int[8]),.T1I1(NET_632),.T1I2(NET_508),.T1I3(p3_fsm[2]),.TB1S(GND),.Q1Z(m1_oper1_raddr_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_Z31_2 (.tFragBitInfo(16'b0111111110000000),.bFragBitInfo(16'b1000000000000000),.B2I0(m1_oper1_raddr_dup_0[7]),.B2I1(m1_oper1_raddr_dup_0[6]),.B2I2(m1_oper1_raddr_dup_0[8]),.B2I3(NET_572),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_raddr_dup_0[3]),.T2I1(m1_oper1_raddr_dup_0[2]),.T2I2(m1_oper1_raddr_dup_0[4]),.T2I3(m1_oper1_raddr_dup_0[5]),.TB2S(GND),.B2Z(NET_652),.C2Z(NET_550),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_Z31_3 (.tFragBitInfo(16'b1110001011000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36808z2),.QCK(CLK_int_0__CAND0_BRSBR_26_padClk),.QRT(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF),.QST(GND),.T3I0(NET_550),.T3I1(NET_508),.T3I2(lint_ADDR_int[5]),.T3I3(p3_fsm[2]),.TB3S(GND),.Q3Z(m1_oper1_raddr_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AA5_0 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx36058z2_CAND4_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(nx11312z1_CAND3_TRSTR_27_tpGCLKBUF),.T0I1(lint_WDATA_int[15]),.T0I2(GND),.T0I3(m0_oper1_rdata_int[15]),.TB0S(GND),.Q0Z(tcdm_wdata_p1_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA5_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA6_0 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx36058z2_CAND4_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(nx11312z1_CAND3_TRSTR_27_tpGCLKBUF),.T0I1(GND),.T0I2(lint_WDATA_int[16]),.T0I3(m0_oper1_rdata_int[16]),.TB0S(GND),.Q0Z(tcdm_wdata_p1_dup_0[16]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA6_1 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx36058z2_CAND4_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T1I0(nx11312z1_CAND3_TRSTR_27_tpGCLKBUF),.T1I1(m0_oper1_rdata_int[18]),.T1I2(lint_WDATA_int[18]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p1_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA6_2 (.tFragBitInfo(16'b0000111000000100),.bFragBitInfo(16'b0111100011110000),.B2I0(tcdm_addr_p0_dup_0[2]),.B2I1(tcdm_addr_p0_dup_0[3]),.B2I2(tcdm_addr_p0_dup_0[5]),.B2I3(tcdm_addr_p0_dup_0[4]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T2I0(nx45272z2),.T2I1(NET_693),.T2I2(GND),.T2I3(lint_WDATA_int[5]),.TB2S(GND),.B2Z(NET_693),.Q2Z(tcdm_addr_p0_dup_0[5]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA6_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36058z2_CAND4_TRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[17]),.T3I1(m0_oper1_rdata_int[17]),.T3I2(nx11312z1_CAND3_TRSTR_27_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p1_dup_0[17]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AA7_0 (.tFragBitInfo(16'b1111011000000110),.bFragBitInfo(16'b0111111110000000),.B0I0(tcdm_addr_p0_dup_0[13]),.B0I1(NET_788),.B0I2(tcdm_addr_p0_dup_0[12]),.B0I3(tcdm_addr_p0_dup_0[14]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(tcdm_addr_p0_dup_0[6]),.T0I1(NET_716),.T0I2(nx45272z2),.T0I3(lint_WDATA_int[6]),.TB0S(GND),.B0Z(NET_787),.Q0Z(tcdm_addr_p0_dup_0[6]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA7_1 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T1I0(nx45272z2),.T1I1(lint_WDATA_int[14]),.T1I2(NET_787),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_addr_p0_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(tcdm_addr_p0_dup_0[4]),.B2I1(tcdm_addr_p0_dup_0[5]),.B2I2(tcdm_addr_p0_dup_0[3]),.B2I3(tcdm_addr_p0_dup_0[2]),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.B2Z(NET_716),.B2CO(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA7_3 (.tFragBitInfo(16'b1011111000010100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T3I0(nx45272z2),.T3I1(NET_788),.T3I2(tcdm_addr_p0_dup_0[12]),.T3I3(lint_WDATA_int[12]),.TB3S(GND),.Q3Z(tcdm_addr_p0_dup_0[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AA8_0 (.tFragBitInfo(16'b1100110001011010),.bFragBitInfo(16'b0111111110000000),.B0I0(tcdm_addr_p0_dup_0[6]),.B0I1(tcdm_addr_p0_dup_0[7]),.B0I2(NET_716),.B0I3(tcdm_addr_p0_dup_0[8]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(tcdm_addr_p0_dup_0[10]),.T0I1(lint_WDATA_int[10]),.T0I2(NET_715),.T0I3(nx45272z2),.TB0S(GND),.B0Z(NET_743),.Q0Z(tcdm_addr_p0_dup_0[10]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA8_1 (.tFragBitInfo(16'b0001010101000000),.bFragBitInfo(16'b1111011011111100),.B1I0(NET_716),.B1I1(tcdm_addr_p0_dup_0[7]),.B1I2(nx45272z2),.B1I3(tcdm_addr_p0_dup_0[6]),.CD1S(GND),.Q1DI(GND),.Q1EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T1I0(nx45272z2),.T1I1(tcdm_addr_p0_dup_0[6]),.T1I2(NET_716),.T1I3(tcdm_addr_p0_dup_0[7]),.TB1S(lint_WDATA_int[7]),.Q1Z(tcdm_addr_p0_dup_0[7]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA8_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B2I0(tcdm_addr_p0_dup_0[6]),.B2I1(tcdm_addr_p0_dup_0[7]),.B2I2(NET_716),.B2I3(tcdm_addr_p0_dup_0[8]),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p0_dup_0[6]),.T2I1(tcdm_addr_p0_dup_0[7]),.T2I2(NET_716),.T2I3(tcdm_addr_p0_dup_0[8]),.TB2S(tcdm_addr_p0_dup_0[9]),.C2Z(NET_715),.B2CO(),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_AA8_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSTR_27_padClk),.QRT(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[8]),.T3I1(NET_743),.T3I2(nx45272z2),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_addr_p0_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AA9_0 (.tFragBitInfo(16'b1100010111001010),.bFragBitInfo(16'b0010000000000000),.B0I0(tcdm_addr_p0_dup_0[13]),.B0I1(GND),.B0I2(tcdm_addr_p0_dup_0[15]),.B0I3(tcdm_addr_p0_dup_0[14]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T0I0(NET_713),.T0I1(lint_WDATA_int[13]),.T0I2(nx45272z2),.T0I3(tcdm_addr_p0_dup_0[13]),.TB0S(GND),.B0Z(NET_714),.Q0Z(tcdm_addr_p0_dup_0[13]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B1I0(NET_714),.B1I1(tcdm_addr_p0_dup_0[16]),.B1I2(NET_713),.B1I3(tcdm_addr_p0_dup_0[17]),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T1I0(NET_713),.T1I1(tcdm_addr_p0_dup_0[17]),.T1I2(NET_714),.T1I3(tcdm_addr_p0_dup_0[16]),.TB1S(tcdm_addr_p0_dup_0[18]),.C1Z(NET_712),.B1CO(),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_AA9_2 (.tFragBitInfo(16'b1010101000111100),.bFragBitInfo(16'b1000000000000000),.B2I0(NET_715),.B2I1(tcdm_addr_p0_dup_0[12]),.B2I2(tcdm_addr_p0_dup_0[10]),.B2I3(tcdm_addr_p0_dup_0[11]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[19]),.T2I1(tcdm_addr_p0_dup_0[19]),.T2I2(NET_712),.T2I3(nx45272z2),.TB2S(GND),.B2Z(NET_713),.Q2Z(tcdm_addr_p0_dup_0[19]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA9_3 (.tFragBitInfo(16'b0000011100001000),.bFragBitInfo(16'b1011111011101110),.B3I0(nx45272z2),.B3I1(tcdm_addr_p0_dup_0[16]),.B3I2(NET_713),.B3I3(NET_714),.CD3S(GND),.Q3DI(GND),.Q3EN(nx42281z2),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T3I0(NET_713),.T3I1(NET_714),.T3I2(nx45272z2),.T3I3(tcdm_addr_p0_dup_0[16]),.TB3S(lint_WDATA_int[16]),.Q3Z(tcdm_addr_p0_dup_0[16]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AA10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.CD0S(VCC),.Q0DI(lint_WDATA_int[0]),.Q0EN(nx45272z2),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.Q0Z(tcdm_addr_p0_dup_0[0]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA10_2 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx36058z2_CAND5_TRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[13]),.T2I1(GND),.T2I2(nx11312z1_CAND4_TRSBR_27_tpGCLKBUF),.T2I3(m0_oper1_rdata_int[13]),.TB2S(GND),.Q2Z(tcdm_wdata_p1_dup_0[13]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA11_0 (.tFragBitInfo(16'b1010001110101100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx13970z2_CAND2_TRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[6]),.T0I1(tcdm_addr_p1_dup_0[6]),.T0I2(nx12973z2_CAND3_TRSBR_27_tpGCLKBUF),.T0I3(NET_330),.TB0S(GND),.Q0Z(tcdm_addr_p1_dup_0[6]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA11_1 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx36058z2_CAND5_TRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T1I0(nx11312z1_CAND4_TRSBR_27_tpGCLKBUF),.T1I1(lint_WDATA_int[14]),.T1I2(m0_oper1_rdata_int[14]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p1_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA11_2 (.tFragBitInfo(16'b0001001000110000),.bFragBitInfo(16'b1101111011111100),.B2I0(tcdm_addr_p1_dup_0[6]),.B2I1(NET_89),.B2I2(tcdm_addr_p1_dup_0[7]),.B2I3(NET_330),.CD2S(GND),.Q2DI(GND),.Q2EN(nx13970z2_CAND2_TRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p1_dup_0[6]),.T2I1(NET_89),.T2I2(tcdm_addr_p1_dup_0[7]),.T2I3(NET_330),.TB2S(lint_WDATA_int[7]),.Q2Z(tcdm_addr_p1_dup_0[7]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA11_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T3I0(tcdm_addr_p1_dup_0[5]),.T3I1(tcdm_addr_p1_dup_0[3]),.T3I2(tcdm_addr_p1_dup_0[4]),.T3I3(tcdm_addr_p1_dup_0[2]),.TB3S(GND),.C3Z(NET_330),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_AA12_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_329),.B0I1(tcdm_addr_p1_dup_0[13]),.B0I2(NET_328),.B0I3(tcdm_addr_p1_dup_0[14]),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T0I0(NET_329),.T0I1(tcdm_addr_p1_dup_0[13]),.T0I2(NET_328),.T0I3(tcdm_addr_p1_dup_0[14]),.TB0S(tcdm_addr_p1_dup_0[15]),.C0Z(NET_327),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA12_1 (.tFragBitInfo(16'b1101111000010010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx13970z2_CAND2_TRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T1I0(NET_459),.T1I1(nx12973z2_CAND3_TRSBR_27_tpGCLKBUF),.T1I2(tcdm_addr_p1_dup_0[13]),.T1I3(lint_WDATA_int[13]),.TB1S(GND),.Q1Z(tcdm_addr_p1_dup_0[13]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA12_2 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'b0000000000100000),.B2I0(NET_329),.B2I1(GND),.B2I2(NET_328),.B2I3(GND),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p1_dup_0[12]),.T2I1(tcdm_addr_p1_dup_0[9]),.T2I2(tcdm_addr_p1_dup_0[11]),.T2I3(tcdm_addr_p1_dup_0[10]),.TB2S(GND),.B2Z(NET_459),.C2Z(NET_329),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_AA12_3 (.tFragBitInfo(16'b0001001100100000),.bFragBitInfo(16'b1111111101101100),.B3I0(tcdm_addr_p1_dup_0[13]),.B3I1(tcdm_addr_p1_dup_0[14]),.B3I2(NET_459),.B3I3(NET_89),.CD3S(GND),.Q3DI(GND),.Q3EN(nx13970z2_CAND2_TRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T3I0(NET_459),.T3I1(NET_89),.T3I2(tcdm_addr_p1_dup_0[13]),.T3I3(tcdm_addr_p1_dup_0[14]),.TB3S(lint_WDATA_int[14]),.Q3Z(tcdm_addr_p1_dup_0[14]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AA13_0 (.tFragBitInfo(16'b1011000111100100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx13970z2_CAND2_TRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T0I0(nx12973z2_CAND3_TRSBR_27_tpGCLKBUF),.T0I1(tcdm_addr_p1_dup_0[9]),.T0I2(lint_WDATA_int[9]),.T0I3(NET_328),.TB0S(GND),.Q0Z(tcdm_addr_p1_dup_0[9]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA13_1 (.tFragBitInfo(16'b0000000010000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(VCC),.Q1DI(lint_WDATA_int[0]),.Q1EN(nx12973z2_CAND3_TRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p1_dup_0[12]),.T1I1(tcdm_addr_p1_dup_0[13]),.T1I2(tcdm_addr_p1_dup_0[14]),.T1I3(GND),.TB1S(GND),.C1Z(NET_352),.Q1Z(tcdm_addr_p1_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.T1CO());

	LOGIC_2 QL_INST_AA13_2 (.tFragBitInfo(16'b1100110001011010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx13970z2_CAND2_TRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p1_dup_0[2]),.T2I1(lint_WDATA_int[3]),.T2I2(tcdm_addr_p1_dup_0[3]),.T2I3(nx12973z2_CAND3_TRSBR_27_tpGCLKBUF),.TB2S(GND),.Q2Z(tcdm_addr_p1_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA13_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_27_padClk),.QRT(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF),.QST(GND),.T3I0(tcdm_addr_p1_dup_0[10]),.T3I1(tcdm_addr_p1_dup_0[9]),.T3I2(tcdm_addr_p1_dup_0[11]),.T3I3(NET_328),.TB3S(GND),.C3Z(NET_351),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_AA16_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCK(GND),.QCKS(GND),.QRT(GND),.QST(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA16_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.QCK(GND),.QRT(GND),.QST(GND),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA16_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0000000000000000),.T2I0(NET_50),.T2I1(tcdm_addr_p2_dup_0[9]),.T2I2(NET_253),.T2I3(tcdm_addr_p1_dup_0[9]),.TB2S(GND),.C2Z(NET_249),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.QCK(GND),.QRT(GND),.QST(GND),.T2CO());

	LOGIC_3 QL_INST_AA16_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.QCK(GND),.QRT(GND),.QST(GND),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA17_0 (.tFragBitInfo(16'b1010001110101100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[3]),.T0I1(tcdm_addr_p2_dup_0[3]),.T0I2(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.T0I3(tcdm_addr_p2_dup_0[2]),.TB0S(GND),.Q0Z(tcdm_addr_p2_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA17_1 (.tFragBitInfo(16'b0000011101110111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T1I0(NET_50),.T1I1(tcdm_addr_p1_dup_0[10]),.T1I2(tcdm_addr_p2_dup_0[10]),.T1I3(NET_253),.C1Z(NET_278),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_AA17_2 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'b0001001101011111),.B2I0(NET_50),.B2I1(tcdm_addr_p2_dup_0[8]),.B2I2(tcdm_addr_p1_dup_0[8]),.B2I3(NET_253),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p2_dup_0[14]),.T2I1(NET_50),.T2I2(tcdm_addr_p1_dup_0[14]),.T2I3(NET_253),.TB2S(GND),.B2Z(NET_386),.C2Z(NET_358),.B2CO(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_AA17_3 (.tFragBitInfo(16'b0001010100111111),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T3I0(NET_50),.T3I1(tcdm_addr_p2_dup_0[3]),.T3I2(NET_253),.T3I3(tcdm_addr_p1_dup_0[3]),.C3Z(NET_888),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_AA18_0 (.tFragBitInfo(16'b0000111000000100),.bFragBitInfo(16'b1000000000000000),.B0I0(tcdm_addr_p2_dup_0[8]),.B0I1(tcdm_addr_p2_dup_0[7]),.B0I2(NET_205),.B0I3(tcdm_addr_p2_dup_0[6]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.T0I1(NET_674),.T0I2(GND),.T0I3(lint_WDATA_int[11]),.TB0S(GND),.B0Z(NET_256),.Q0Z(tcdm_addr_p2_dup_0[11]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA18_1 (.tFragBitInfo(16'b0001010001000100),.bFragBitInfo(16'b1111011111111000),.B1I0(NET_205),.B1I1(tcdm_addr_p2_dup_0[6]),.B1I2(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.B1I3(tcdm_addr_p2_dup_0[7]),.CD1S(GND),.Q1DI(GND),.Q1EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T1I0(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.T1I1(tcdm_addr_p2_dup_0[7]),.T1I2(NET_205),.T1I3(tcdm_addr_p2_dup_0[6]),.TB1S(lint_WDATA_int[7]),.Q1Z(tcdm_addr_p2_dup_0[7]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA18_2 (.tFragBitInfo(16'b0110101010101010),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p2_dup_0[11]),.T2I1(NET_256),.T2I2(tcdm_addr_p2_dup_0[9]),.T2I3(tcdm_addr_p2_dup_0[10]),.TB2S(GND),.C2Z(NET_674),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO());

	LOGIC_3 QL_INST_AA18_3 (.tFragBitInfo(16'b1010001110101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[9]),.T3I1(NET_256),.T3I2(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.T3I3(tcdm_addr_p2_dup_0[9]),.TB3S(GND),.Q3Z(tcdm_addr_p2_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AA19_0 (.tFragBitInfo(16'b0101000001000100),.bFragBitInfo(16'b0110101010101010),.B0I0(tcdm_addr_p2_dup_0[15]),.B0I1(NET_717),.B0I2(tcdm_addr_p2_dup_0[13]),.B0I3(tcdm_addr_p2_dup_0[14]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(NET_746),.T0I2(lint_WDATA_int[15]),.T0I3(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.TB0S(GND),.B0Z(NET_746),.Q0Z(tcdm_addr_p2_dup_0[15]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA19_1 (.tFragBitInfo(16'b0000011100001000),.bFragBitInfo(16'b1011111011101110),.B1I0(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.B1I1(tcdm_addr_p2_dup_0[14]),.B1I2(NET_717),.B1I3(tcdm_addr_p2_dup_0[13]),.CD1S(GND),.Q1DI(GND),.Q1EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T1I0(NET_717),.T1I1(tcdm_addr_p2_dup_0[13]),.T1I2(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.T1I3(tcdm_addr_p2_dup_0[14]),.TB1S(lint_WDATA_int[14]),.Q1Z(tcdm_addr_p2_dup_0[14]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA19_2 (.tFragBitInfo(16'b1111000001100110),.bFragBitInfo(16'b0000100000000000),.B2I0(tcdm_addr_p2_dup_0[15]),.B2I1(tcdm_addr_p2_dup_0[13]),.B2I2(GND),.B2I3(tcdm_addr_p2_dup_0[14]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p2_dup_0[13]),.T2I1(NET_717),.T2I2(lint_WDATA_int[13]),.T2I3(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.TB2S(GND),.B2Z(NET_765),.Q2Z(tcdm_addr_p2_dup_0[13]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA19_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B3I0(tcdm_addr_p2_dup_0[11]),.B3I1(tcdm_addr_p2_dup_0[10]),.B3I2(NET_765),.B3I3(NET_651),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T3I0(NET_765),.T3I1(NET_651),.T3I2(tcdm_addr_p2_dup_0[11]),.T3I3(tcdm_addr_p2_dup_0[10]),.TB3S(tcdm_addr_p2_dup_0[12]),.C3Z(NET_764),.B3CO(),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO());

	LOGIC_0 QL_INST_AA20_0 (.tFragBitInfo(16'b1111000001100110),.bFragBitInfo(16'b1000000000000000),.B0I0(tcdm_addr_p2_dup_0[16]),.B0I1(NET_764),.B0I2(tcdm_addr_p2_dup_0[17]),.B0I3(tcdm_addr_p2_dup_0[18]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(tcdm_addr_p2_dup_0[16]),.T0I1(NET_764),.T0I2(lint_WDATA_int[16]),.T0I3(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.TB0S(GND),.B0Z(NET_814),.Q0Z(tcdm_addr_p2_dup_0[16]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA20_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T1I0(NET_812),.T1I1(lint_WDATA_int[18]),.T1I2(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_addr_p2_dup_0[18]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA20_2 (.tFragBitInfo(16'b1111000001100110),.bFragBitInfo(16'b0111111110000000),.B2I0(tcdm_addr_p2_dup_0[16]),.B2I1(NET_764),.B2I2(tcdm_addr_p2_dup_0[17]),.B2I3(tcdm_addr_p2_dup_0[18]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p2_dup_0[19]),.T2I1(NET_814),.T2I2(lint_WDATA_int[19]),.T2I3(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.TB2S(GND),.B2Z(NET_812),.Q2Z(tcdm_addr_p2_dup_0[19]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA20_3 (.tFragBitInfo(16'b0000011100001000),.bFragBitInfo(16'b1011111011101110),.B3I0(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.B3I1(tcdm_addr_p2_dup_0[17]),.B3I2(tcdm_addr_p2_dup_0[16]),.B3I3(NET_764),.CD3S(GND),.Q3DI(GND),.Q3EN(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T3I0(tcdm_addr_p2_dup_0[16]),.T3I1(NET_764),.T3I2(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF),.T3I3(tcdm_addr_p2_dup_0[17]),.TB3S(lint_WDATA_int[17]),.Q3Z(tcdm_addr_p2_dup_0[17]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AA21_0 (.tFragBitInfo(16'b1010101000111100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60936z2_CAND5_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[15]),.T0I1(tcdm_addr_p3_dup_0[15]),.T0I2(NET_301),.T0I3(nx40548z2_CAND3_BRSTR_27_tpGCLKBUF),.TB0S(GND),.Q0Z(tcdm_addr_p3_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA21_1 (.tFragBitInfo(16'b0001001000110000),.bFragBitInfo(16'b1111111101101010),.B1I0(tcdm_addr_p3_dup_0[19]),.B1I1(NET_845),.B1I2(tcdm_addr_p3_dup_0[15]),.B1I3(nx40548z2_CAND3_BRSTR_27_tpGCLKBUF),.CD1S(GND),.Q1DI(GND),.Q1EN(nx60936z2_CAND5_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p3_dup_0[15]),.T1I1(nx40548z2_CAND3_BRSTR_27_tpGCLKBUF),.T1I2(tcdm_addr_p3_dup_0[19]),.T1I3(NET_845),.TB1S(lint_WDATA_int[19]),.Q1Z(tcdm_addr_p3_dup_0[19]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA21_2 (.tFragBitInfo(16'b0000000001101100),.bFragBitInfo(16'b1111111101101100),.B2I0(tcdm_addr_p3_dup_0[15]),.B2I1(tcdm_addr_p3_dup_0[16]),.B2I2(NET_301),.B2I3(nx40548z2_CAND3_BRSTR_27_tpGCLKBUF),.CD2S(GND),.Q2DI(GND),.Q2EN(nx60936z2_CAND5_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p3_dup_0[15]),.T2I1(tcdm_addr_p3_dup_0[16]),.T2I2(NET_301),.T2I3(nx40548z2_CAND3_BRSTR_27_tpGCLKBUF),.TB2S(lint_WDATA_int[16]),.Q2Z(tcdm_addr_p3_dup_0[16]),.B2CO(),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA21_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T3I0(tcdm_addr_p3_dup_0[18]),.T3I1(tcdm_addr_p3_dup_0[16]),.T3I2(tcdm_addr_p3_dup_0[17]),.T3I3(NET_301),.C3Z(NET_845),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_AA22_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AA22_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AA22_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AA22_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(tcdm_rdata_p3_int[15]),.Q3EN(tcdm_valid_p3_int),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.Q3Z(tcdm_result_p3[15]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA23_0 (.tFragBitInfo(16'b0100010001010000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60936z2_CAND5_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(lint_WDATA_int[5]),.T0I2(NET_820),.T0I3(nx40548z2_CAND3_BRSTR_27_tpGCLKBUF),.TB0S(GND),.Q0Z(tcdm_addr_p3_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA23_1 (.tFragBitInfo(16'b0111111110000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p3_dup_0[2]),.T1I1(tcdm_addr_p3_dup_0[3]),.T1I2(tcdm_addr_p3_dup_0[4]),.T1I3(tcdm_addr_p3_dup_0[5]),.C1Z(NET_820),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_AA23_2 (.tFragBitInfo(16'b1111000001100110),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx60936z2_CAND5_BRSTR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T2I0(tcdm_addr_p3_dup_0[2]),.T2I1(tcdm_addr_p3_dup_0[3]),.T2I2(lint_WDATA_int[3]),.T2I3(nx40548z2_CAND3_BRSTR_27_tpGCLKBUF),.TB2S(GND),.Q2Z(tcdm_addr_p3_dup_0[3]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA23_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AA24_0 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T0I0(nx3850z2),.T0I1(lint_WDATA_int[3]),.T0I2(GND),.T0I3(tcdm_rdata_p3_int[3]),.TB0S(GND),.Q0Z(m1_oper1_wdata_dup_0[3]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA24_1 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T1I0(nx3850z2),.T1I1(tcdm_rdata_p3_int[5]),.T1I2(lint_WDATA_int[5]),.T1I3(GND),.TB1S(GND),.Q1Z(m1_oper1_wdata_dup_0[5]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA24_2 (.tFragBitInfo(16'b0011001000010000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T2I0(nx3850z2),.T2I1(GND),.T2I2(tcdm_rdata_p3_int[2]),.T2I3(lint_WDATA_int[2]),.TB2S(GND),.Q2Z(m1_oper1_wdata_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA24_3 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx3786z2),.QCK(CLK_int_0__CAND0_BRSTR_27_padClk),.QRT(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF),.QST(GND),.T3I0(nx3850z2),.T3I1(tcdm_rdata_p3_int[7]),.T3I2(lint_WDATA_int[7]),.T3I3(GND),.TB3S(GND),.Q3Z(m1_oper1_wdata_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AA25_0 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx3786z2_CAND5_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND2_BRSBR_27_tpGCLKBUF),.QST(GND),.T0I0(nx3850z2_CAND3_BRSBR_27_tpGCLKBUF),.T0I1(lint_WDATA_int[15]),.T0I2(GND),.T0I3(tcdm_rdata_p3_int[15]),.TB0S(GND),.Q0Z(m1_oper1_wdata_dup_0[15]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA25_1 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx25788z3_CAND4_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND2_BRSBR_27_tpGCLKBUF),.QST(GND),.T1I0(m1_oper1_rdata_int[14]),.T1I1(lint_WDATA_int[14]),.T1I2(NET_0_CAND1_BRSBR_27_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p3_dup_0[14]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA25_2 (.tFragBitInfo(16'b0000110000001010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx25788z3_CAND4_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND2_BRSBR_27_tpGCLKBUF),.QST(GND),.T2I0(m1_oper1_rdata_int[15]),.T2I1(lint_WDATA_int[15]),.T2I2(GND),.T2I3(NET_0_CAND1_BRSBR_27_tpGCLKBUF),.TB2S(GND),.Q2Z(tcdm_wdata_p3_dup_0[15]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA25_3 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx25788z3_CAND4_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND2_BRSBR_27_tpGCLKBUF),.QST(GND),.T3I0(m1_oper1_rdata_int[13]),.T3I1(lint_WDATA_int[13]),.T3I2(NET_0_CAND1_BRSBR_27_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p3_dup_0[13]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AA26_0 (.tFragBitInfo(16'b0000111000000100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx25788z3_CAND4_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND2_BRSBR_27_tpGCLKBUF),.QST(GND),.T0I0(NET_0_CAND1_BRSBR_27_tpGCLKBUF),.T0I1(m1_oper1_rdata_int[18]),.T0I2(GND),.T0I3(lint_WDATA_int[18]),.TB0S(GND),.Q0Z(tcdm_wdata_p3_dup_0[18]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AA26_1 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx25788z3_CAND4_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND2_BRSBR_27_tpGCLKBUF),.QST(GND),.T1I0(NET_0_CAND1_BRSBR_27_tpGCLKBUF),.T1I1(lint_WDATA_int[17]),.T1I2(GND),.T1I3(m1_oper1_rdata_int[17]),.TB1S(GND),.Q1Z(tcdm_wdata_p3_dup_0[17]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AA26_2 (.tFragBitInfo(16'b0000101000001100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx25788z3_CAND4_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND2_BRSBR_27_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[19]),.T2I1(m1_oper1_rdata_int[19]),.T2I2(GND),.T2I3(NET_0_CAND1_BRSBR_27_tpGCLKBUF),.TB2S(GND),.Q2Z(tcdm_wdata_p3_dup_0[19]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AA26_3 (.tFragBitInfo(16'b0010001000110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx25788z3_CAND4_BRSBR_27_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_27_padClk),.QRT(not_RESET_0_CAND2_BRSBR_27_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[16]),.T3I1(GND),.T3I2(m1_oper1_rdata_int[16]),.T3I3(NET_0_CAND1_BRSBR_27_tpGCLKBUF),.TB3S(GND),.Q3Z(tcdm_wdata_p3_dup_0[16]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB4_2 (.tFragBitInfo(16'b0000111000000010),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx36058z2_CAND4_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.T2I0(m0_oper1_rdata_int[7]),.T2I1(nx11312z1_CAND3_TRSTR_28_tpGCLKBUF),.T2I2(GND),.T2I3(lint_WDATA_int[7]),.TB2S(GND),.Q2Z(tcdm_wdata_p1_dup_0[7]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AB4_3 (.tFragBitInfo(16'b0000000011001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36058z2_CAND4_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.T3I0(m0_oper1_rdata_int[6]),.T3I1(lint_WDATA_int[6]),.T3I2(nx11312z1_CAND3_TRSTR_28_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p1_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB6_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB6_1 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx36058z2_CAND4_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.T1I0(m0_oper1_rdata_int[12]),.T1I1(nx11312z1_CAND3_TRSTR_28_tpGCLKBUF),.T1I2(lint_WDATA_int[12]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p1_dup_0[12]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AB6_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB6_3 (.tFragBitInfo(16'b0000000010111000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36058z2_CAND4_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[8]),.T3I1(nx11312z1_CAND3_TRSTR_28_tpGCLKBUF),.T3I2(m0_oper1_rdata_int[8]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p1_dup_0[8]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB7_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB7_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB7_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB7_3 (.tFragBitInfo(16'b0011001000000010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36058z2_CAND4_TRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_28_padClk),.QRT(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF),.QST(GND),.T3I0(m0_oper1_rdata_int[11]),.T3I1(GND),.T3I2(nx11312z1_CAND3_TRSTR_28_tpGCLKBUF),.T3I3(lint_WDATA_int[11]),.TB3S(GND),.Q3Z(tcdm_wdata_p1_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB9_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB9_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36058z2_CAND5_TRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[9]),.T3I1(m0_oper1_rdata_int[9]),.T3I2(nx11312z1_CAND4_TRSBR_28_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p1_dup_0[9]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB10_0 (.tFragBitInfo(16'b0010001100100000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx36058z2_CAND5_TRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.T0I0(lint_WDATA_int[4]),.T0I1(GND),.T0I2(nx11312z1_CAND4_TRSBR_28_tpGCLKBUF),.T0I3(m0_oper1_rdata_int[4]),.TB0S(GND),.Q0Z(tcdm_wdata_p1_dup_0[4]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AB10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB10_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AB11_0 (.tFragBitInfo(16'b0000011000001010),.bFragBitInfo(16'b1111011011111010),.B0I0(tcdm_addr_p1_dup_0[10]),.B0I1(tcdm_addr_p1_dup_0[9]),.B0I2(NET_89),.B0I3(NET_328),.CD0S(GND),.Q0DI(GND),.Q0EN(nx13970z2_CAND2_TRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.T0I0(tcdm_addr_p1_dup_0[10]),.T0I1(tcdm_addr_p1_dup_0[9]),.T0I2(NET_89),.T0I3(NET_328),.TB0S(lint_WDATA_int[10]),.Q0Z(tcdm_addr_p1_dup_0[10]),.B0CO(),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AB11_1 (.tFragBitInfo(16'b0101010000000100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx13970z2_CAND2_TRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.T1I0(GND),.T1I1(NET_868),.T1I2(NET_89),.T1I3(lint_WDATA_int[8]),.TB1S(GND),.Q1Z(tcdm_addr_p1_dup_0[8]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AB11_2 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0111100011110000),.B2I0(NET_330),.B2I1(tcdm_addr_p1_dup_0[6]),.B2I2(tcdm_addr_p1_dup_0[8]),.B2I3(tcdm_addr_p1_dup_0[7]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx36058z2_CAND5_TRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.T2I0(nx11312z1_CAND4_TRSBR_28_tpGCLKBUF),.T2I1(lint_WDATA_int[10]),.T2I2(GND),.T2I3(m0_oper1_rdata_int[10]),.TB2S(GND),.B2Z(NET_868),.Q2Z(tcdm_wdata_p1_dup_0[10]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AB11_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.T3I0(NET_330),.T3I1(tcdm_addr_p1_dup_0[6]),.T3I2(tcdm_addr_p1_dup_0[8]),.T3I3(tcdm_addr_p1_dup_0[7]),.C3Z(NET_328),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.TB3S(GND));

	LOGIC_0 QL_INST_AB12_0 (.tFragBitInfo(16'b0101000001000100),.bFragBitInfo(16'b0110101010101010),.B0I0(tcdm_addr_p1_dup_0[5]),.B0I1(tcdm_addr_p1_dup_0[2]),.B0I2(tcdm_addr_p1_dup_0[3]),.B0I3(tcdm_addr_p1_dup_0[4]),.CD0S(GND),.Q0DI(GND),.Q0EN(nx13970z2_CAND2_TRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.T0I0(GND),.T0I1(NET_88),.T0I2(lint_WDATA_int[5]),.T0I3(NET_89),.TB0S(GND),.B0Z(NET_88),.Q0Z(tcdm_addr_p1_dup_0[5]),.B0CO(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AB12_1 (.tFragBitInfo(16'b0110110011001100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p1_dup_0[9]),.T1I1(tcdm_addr_p1_dup_0[11]),.T1I2(tcdm_addr_p1_dup_0[10]),.T1I3(NET_328),.TB1S(GND),.C1Z(NET_511),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_AB12_2 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx13970z2_CAND2_TRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_WDATA_int[11]),.T2I2(NET_89),.T2I3(NET_511),.TB2S(GND),.Q2Z(tcdm_addr_p1_dup_0[11]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AB12_3 (.tFragBitInfo(16'b0001010101000000),.bFragBitInfo(16'b1111011011111100),.B3I0(tcdm_addr_p1_dup_0[3]),.B3I1(tcdm_addr_p1_dup_0[4]),.B3I2(NET_89),.B3I3(tcdm_addr_p1_dup_0[2]),.CD3S(GND),.Q3DI(GND),.Q3EN(nx13970z2_CAND2_TRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_28_padClk),.QRT(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF),.QST(GND),.T3I0(NET_89),.T3I1(tcdm_addr_p1_dup_0[2]),.T3I2(tcdm_addr_p1_dup_0[3]),.T3I3(tcdm_addr_p1_dup_0[4]),.TB3S(lint_WDATA_int[4]),.Q3Z(tcdm_addr_p1_dup_0[4]),.B3CO(),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB17_0 (.tFragBitInfo(16'b0011000000100010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx60851z2_CAND4_BRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T0I0(NET_848),.T0I1(GND),.T0I2(lint_WDATA_int[5]),.T0I3(nx63842z2_CAND1_BRSTR_28_tpGCLKBUF),.TB0S(GND),.Q0Z(tcdm_addr_p2_dup_0[5]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AB17_1 (.tFragBitInfo(16'b0000011100001000),.bFragBitInfo(16'b1011111011101110),.B1I0(nx63842z2_CAND1_BRSTR_28_tpGCLKBUF),.B1I1(tcdm_addr_p2_dup_0[4]),.B1I2(tcdm_addr_p2_dup_0[2]),.B1I3(tcdm_addr_p2_dup_0[3]),.CD1S(GND),.Q1DI(GND),.Q1EN(nx60851z2_CAND4_BRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p2_dup_0[2]),.T1I1(tcdm_addr_p2_dup_0[3]),.T1I2(nx63842z2_CAND1_BRSTR_28_tpGCLKBUF),.T1I3(tcdm_addr_p2_dup_0[4]),.TB1S(lint_WDATA_int[4]),.Q1Z(tcdm_addr_p2_dup_0[4]),.B1CO(),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AB17_2 (.tFragBitInfo(16'b0000101000000011),.bFragBitInfo(16'b0110101010101010),.B2I0(tcdm_addr_p2_dup_0[5]),.B2I1(tcdm_addr_p2_dup_0[3]),.B2I2(tcdm_addr_p2_dup_0[2]),.B2I3(tcdm_addr_p2_dup_0[4]),.CD2S(GND),.Q2DI(GND),.Q2EN(nx60851z2_CAND4_BRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T2I0(lint_WDATA_int[2]),.T2I1(tcdm_addr_p2_dup_0[2]),.T2I2(GND),.T2I3(nx63842z2_CAND1_BRSTR_28_tpGCLKBUF),.TB2S(GND),.B2Z(NET_848),.Q2Z(tcdm_addr_p2_dup_0[2]),.B2CO(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AB17_3 (.tFragBitInfo(16'b1000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(VCC),.Q3DI(lint_WDATA_int[1]),.Q3EN(nx63842z2_CAND1_BRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T3I0(tcdm_addr_p2_dup_0[5]),.T3I1(tcdm_addr_p2_dup_0[3]),.T3I2(tcdm_addr_p2_dup_0[2]),.T3I3(tcdm_addr_p2_dup_0[4]),.TB3S(GND),.C3Z(NET_205),.Q3Z(tcdm_addr_p2_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.T3CO());

	LOGIC_0 QL_INST_AB18_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(tcdm_addr_p2_dup_0[8]),.B0I1(tcdm_addr_p2_dup_0[7]),.B0I2(tcdm_addr_p2_dup_0[6]),.B0I3(NET_205),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T0I0(tcdm_addr_p2_dup_0[8]),.T0I1(tcdm_addr_p2_dup_0[7]),.T0I2(tcdm_addr_p2_dup_0[6]),.T0I3(NET_205),.TB0S(tcdm_addr_p2_dup_0[9]),.C0Z(NET_651),.B0CO(),.B0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AB18_1 (.tFragBitInfo(16'b0110101010101010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T1I0(tcdm_addr_p2_dup_0[8]),.T1I1(tcdm_addr_p2_dup_0[7]),.T1I2(NET_205),.T1I3(tcdm_addr_p2_dup_0[6]),.TB1S(GND),.C1Z(NET_203),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO());

	LOGIC_2 QL_INST_AB18_2 (.tFragBitInfo(16'b0100010101000000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx60851z2_CAND4_BRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T2I0(GND),.T2I1(lint_WDATA_int[8]),.T2I2(nx63842z2_CAND1_BRSTR_28_tpGCLKBUF),.T2I3(NET_203),.TB2S(GND),.Q2Z(tcdm_addr_p2_dup_0[8]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AB18_3 (.tFragBitInfo(16'b1100010111001010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx60851z2_CAND4_BRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T3I0(NET_205),.T3I1(lint_WDATA_int[6]),.T3I2(nx63842z2_CAND1_BRSTR_28_tpGCLKBUF),.T3I3(tcdm_addr_p2_dup_0[6]),.TB3S(GND),.Q3Z(tcdm_addr_p2_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB19_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b1000000000000000),.B0I0(NET_651),.B0I1(tcdm_addr_p2_dup_0[10]),.B0I2(tcdm_addr_p2_dup_0[11]),.B0I3(tcdm_addr_p2_dup_0[12]),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.B0Z(NET_717),.B0CO(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AB19_1 (.tFragBitInfo(16'b0111100011110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T1I0(NET_651),.T1I1(tcdm_addr_p2_dup_0[10]),.T1I2(tcdm_addr_p2_dup_0[12]),.T1I3(tcdm_addr_p2_dup_0[11]),.C1Z(NET_694),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.TB1S(GND));

	LOGIC_2 QL_INST_AB19_2 (.tFragBitInfo(16'b1111000001100110),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx60851z2_CAND4_BRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T2I0(NET_651),.T2I1(tcdm_addr_p2_dup_0[10]),.T2I2(lint_WDATA_int[10]),.T2I3(nx63842z2_CAND1_BRSTR_28_tpGCLKBUF),.TB2S(GND),.Q2Z(tcdm_addr_p2_dup_0[10]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AB19_3 (.tFragBitInfo(16'b0000000011011000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx60851z2_CAND4_BRSTR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T3I0(nx63842z2_CAND1_BRSTR_28_tpGCLKBUF),.T3I1(lint_WDATA_int[12]),.T3I2(NET_694),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_addr_p2_dup_0[12]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB24_0 (.tFragBitInfo(16'b0000111000000010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx25788z3),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_rdata_int[10]),.T0I1(NET_0),.T0I2(GND),.T0I3(lint_WDATA_int[10]),.TB0S(GND),.Q0Z(tcdm_wdata_p3_dup_0[10]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AB24_1 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx25788z3),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T1I0(NET_0),.T1I1(m1_oper1_rdata_int[4]),.T1I2(lint_WDATA_int[4]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p3_dup_0[4]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AB24_2 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx25788z3),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T2I0(NET_0),.T2I1(m1_oper1_rdata_int[9]),.T2I2(lint_WDATA_int[9]),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_wdata_p3_dup_0[9]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AB24_3 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx25788z3),.QCK(CLK_int_0__CAND0_BRSTR_28_padClk),.QRT(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF),.QST(GND),.T3I0(NET_0),.T3I1(m1_oper1_rdata_int[7]),.T3I2(lint_WDATA_int[7]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p3_dup_0[7]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB25_0 (.tFragBitInfo(16'b0000111000000100),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx25788z3_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND2_BRSBR_28_tpGCLKBUF),.QST(GND),.T0I0(NET_0_CAND1_BRSBR_28_tpGCLKBUF),.T0I1(m1_oper1_rdata_int[8]),.T0I2(GND),.T0I3(lint_WDATA_int[8]),.TB0S(GND),.Q0Z(tcdm_wdata_p3_dup_0[8]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AB25_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND2_BRSBR_28_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB25_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND2_BRSBR_28_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB25_3 (.tFragBitInfo(16'b0010001000110000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx25788z3_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND2_BRSBR_28_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[11]),.T3I1(GND),.T3I2(m1_oper1_rdata_int[11]),.T3I3(NET_0_CAND1_BRSBR_28_tpGCLKBUF),.TB3S(GND),.Q3Z(tcdm_wdata_p3_dup_0[11]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AB26_0 (.tFragBitInfo(16'b0000110100001000),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx25788z3_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND2_BRSBR_28_tpGCLKBUF),.QST(GND),.T0I0(NET_0_CAND1_BRSBR_28_tpGCLKBUF),.T0I1(lint_WDATA_int[12]),.T0I2(GND),.T0I3(m1_oper1_rdata_int[12]),.TB0S(GND),.Q0Z(tcdm_wdata_p3_dup_0[12]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AB26_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND2_BRSBR_28_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AB26_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND2_BRSBR_28_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AB26_3 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx25788z3_CAND4_BRSBR_28_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_28_padClk),.QRT(not_RESET_0_CAND2_BRSBR_28_tpGCLKBUF),.QST(GND),.T3I0(NET_0_CAND1_BRSBR_28_tpGCLKBUF),.T3I1(m1_oper1_rdata_int[6]),.T3I2(lint_WDATA_int[6]),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p3_dup_0[6]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AC4_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC4_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC4_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC4_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36058z2_CAND4_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[0]),.T3I1(m0_oper1_rdata_int[0]),.T3I2(nx11312z1_CAND3_TRSTR_29_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p1_dup_0[0]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AC5_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC5_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC5_2 (.tFragBitInfo(16'b0011000100100000),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx36058z2_CAND4_TRSTR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.T2I0(nx11312z1_CAND3_TRSTR_29_tpGCLKBUF),.T2I1(GND),.T2I2(lint_WDATA_int[2]),.T2I3(m0_oper1_rdata_int[2]),.TB2S(GND),.Q2Z(tcdm_wdata_p1_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AC5_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSTR_29_padClk),.QRT(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	LOGIC_0 QL_INST_AC9_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC9_1 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx36058z2_CAND5_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.T1I0(lint_WDATA_int[3]),.T1I1(m0_oper1_rdata_int[3]),.T1I2(nx11312z1_CAND4_TRSBR_29_tpGCLKBUF),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p1_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AC9_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC9_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36058z2_CAND5_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[1]),.T3I1(m0_oper1_rdata_int[1]),.T3I2(nx11312z1_CAND4_TRSBR_29_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p1_dup_0[1]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AC10_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC10_1 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.CD1S(VCC),.Q1DI(GND),.Q1EN(GND),.Q1Z(),.T1CO(),.T1I0(GND),.T1I1(GND),.T1I2(GND),.T1I3(GND),.TB1S(GND));

	LOGIC_2 QL_INST_AC10_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC10_3 (.tFragBitInfo(16'b0000000010101100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx36058z2_CAND5_TRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_TRSBR_29_padClk),.QRT(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF),.QST(GND),.T3I0(lint_WDATA_int[5]),.T3I1(m0_oper1_rdata_int[5]),.T3I2(nx11312z1_CAND4_TRSBR_29_tpGCLKBUF),.T3I3(GND),.TB3S(GND),.Q3Z(tcdm_wdata_p1_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AC24_0 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'b0000000000000000),.CD0S(GND),.Q0DI(GND),.Q0EN(nx25788z3),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND2_BRSTR_29_tpGCLKBUF),.QST(GND),.T0I0(m1_oper1_rdata_int[1]),.T0I1(NET_0),.T0I2(lint_WDATA_int[1]),.T0I3(GND),.TB0S(GND),.Q0Z(tcdm_wdata_p3_dup_0[1]),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.QCKS(GND),.T0CO());

	LOGIC_1 QL_INST_AC24_1 (.tFragBitInfo(16'b0000000011100010),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx25788z3),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND2_BRSTR_29_tpGCLKBUF),.QST(GND),.T1I0(m1_oper1_rdata_int[3]),.T1I1(NET_0),.T1I2(lint_WDATA_int[3]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p3_dup_0[3]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AC24_2 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND2_BRSTR_29_tpGCLKBUF),.QST(GND),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.CD2S(VCC),.Q2DI(GND),.Q2EN(GND),.Q2Z(),.T2CO(),.T2I0(GND),.T2I1(GND),.T2I2(GND),.T2I3(GND),.TB2S(GND));

	LOGIC_3 QL_INST_AC24_3 (.tFragBitInfo(16'b0101010000010000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD3S(GND),.Q3DI(GND),.Q3EN(nx25788z3),.QCK(CLK_int_0__CAND0_BRSTR_29_padClk),.QRT(not_RESET_0_CAND2_BRSTR_29_tpGCLKBUF),.QST(GND),.T3I0(GND),.T3I1(NET_0),.T3I2(m1_oper1_rdata_int[5]),.T3I3(lint_WDATA_int[5]),.TB3S(GND),.Q3Z(tcdm_wdata_p3_dup_0[5]),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.T3CO());

	LOGIC_0 QL_INST_AC25_0 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'b0000000000000000),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND2_BRSBR_29_tpGCLKBUF),.QST(GND),.B0CO(),.B0I0(GND),.B0I1(GND),.B0I2(GND),.B0I3(GND),.B0Z(),.C0Z(),.CD0S(VCC),.Q0DI(GND),.Q0EN(GND),.Q0Z(),.QCKS(GND),.T0CO(),.T0I0(GND),.T0I1(GND),.T0I2(GND),.T0I3(GND),.TB0S(GND));

	LOGIC_1 QL_INST_AC25_1 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.CD1S(GND),.Q1DI(GND),.Q1EN(nx25788z3_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND2_BRSBR_29_tpGCLKBUF),.QST(GND),.T1I0(NET_0_CAND1_BRSBR_29_tpGCLKBUF),.T1I1(m1_oper1_rdata_int[0]),.T1I2(lint_WDATA_int[0]),.T1I3(GND),.TB1S(GND),.Q1Z(tcdm_wdata_p3_dup_0[0]),.B1CO(),.B1I0(GND),.B1I1(GND),.B1I2(GND),.B1I3(GND),.B1Z(),.C1Z(),.T1CO());

	LOGIC_2 QL_INST_AC25_2 (.tFragBitInfo(16'b0000000011100100),.bFragBitInfo(16'b0000000000000000),.CD2S(GND),.Q2DI(GND),.Q2EN(nx25788z3_CAND4_BRSBR_29_tpGCLKBUF),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND2_BRSBR_29_tpGCLKBUF),.QST(GND),.T2I0(NET_0_CAND1_BRSBR_29_tpGCLKBUF),.T2I1(m1_oper1_rdata_int[2]),.T2I2(lint_WDATA_int[2]),.T2I3(GND),.TB2S(GND),.Q2Z(tcdm_wdata_p3_dup_0[2]),.B2CO(),.B2I0(GND),.B2I1(GND),.B2I2(GND),.B2I3(GND),.B2Z(),.C2Z(),.T2CO());

	LOGIC_3 QL_INST_AC25_3 (.tFragBitInfo(16'b0000000000000000),.bFragBitInfo(16'bxxxxxxxxxxxxxxxx),.QCK(CLK_int_0__CAND0_BRSBR_29_padClk),.QRT(not_RESET_0_CAND2_BRSBR_29_tpGCLKBUF),.QST(GND),.B3CO(),.B3I0(GND),.B3I1(GND),.B3I2(GND),.B3I3(GND),.B3Z(),.C3Z(),.CD3S(VCC),.Q3DI(GND),.Q3EN(GND),.Q3Z(),.T3CO(),.T3I0(GND),.T3I1(GND),.T3I2(GND),.T3I3(GND),.TB3S(GND));

	CLOCK QL_INST_IO_CLK0 (.CEN(VCC),.IP(CLK[0]),.IC(CLK_int[0]),.OP());

	CLOCK QL_INST_IO_CLK1 (.CEN(VCC),.IP(CLK[1]),.IC(CLK_int[1]),.OP());

	CLOCK QL_INST_IO_CLK2 (.CEN(VCC),.IP(CLK[2]),.IC(CLK_int[2]),.OP());

	CLOCK QL_INST_IO_CLK3 (.CEN(VCC),.IP(CLK[3]),.IC(CLK_int[3]),.OP());

	CLOCK QL_INST_IO_CLK4 (.CEN(VCC),.IP(CLK[4]),.IC(CLK_int[4]),.OP());

	CLOCK QL_INST_IO_CLK5 (.CEN(VCC),.IP(CLK[5]),.IC(CLK_int[5]),.OP());

	GMUX QL_INST_GMUX_0 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[0]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_0__GMUX_0_padClk));

	GMUX QL_INST_GMUX_1 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[1]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_1__GMUX_1_padClk));

	GMUX QL_INST_GMUX_2 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[2]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_2__GMUX_2_padClk));

	GMUX QL_INST_GMUX_3 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[3]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_3__GMUX_3_padClk));

	GMUX QL_INST_GMUX_4 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[4]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_4__GMUX_4_padClk));

	GMUX QL_INST_GMUX_5 (.BL_DEN(GND),.BL_DYNEN(GND),.BL_SEN(VCC),.BL_VLP(GND),.BR_DEN(GND),.BR_DYNEN(GND),.BR_SEN(VCC),.BR_VLP(GND),.GCLKIN(CLK_int[5]),.GHSCK(GND),.SSEL(GND),.TL_DEN(GND),.TL_DYNEN(GND),.TL_SEN(VCC),.TL_VLP(GND),.TR_DEN(GND),.TR_DYNEN(GND),.TR_SEN(VCC),.TR_VLP(GND),.IZ(CLK_int_5__GMUX_5_padClk));

	QPMUX QL_INST_QMUX_TL0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_TL0_padClk));

	QPMUX QL_INST_QMUX_TL1 (.GMUXIN(GND),.IS0(VCC),.IS1(VCC),.QCLKIN(GND),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_TL1_tpGCLKBUF));

	QPMUX QL_INST_QMUX_TR0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_TR0_padClk));

	QPMUX QL_INST_QMUX_TR1 (.GMUXIN(GND),.IS0(VCC),.IS1(VCC),.QCLKIN(GND),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_TR1_tpGCLKBUF));

	QPMUX QL_INST_QMUX_TR2 (.GMUXIN(CLK_int_2__GMUX_2_padClk),.IS0(VCC),.IS1(GND),.QCLKIN(GND),.QHSCK(GND),.IZ(CLK_int_2__QMUX_TR2_padClk));

	QMUX QL_INST_QMUX_TR3 (.GMUXIN(CLK_int_3__GMUX_3_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_3__QMUX_TR3_padClk));

	QMUX QL_INST_QMUX_TR4 (.GMUXIN(CLK_int_4__GMUX_4_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_4__QMUX_TR4_padClk));

	QMUX QL_INST_QMUX_TR5 (.GMUXIN(CLK_int_5__GMUX_5_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_5__QMUX_TR5_padClk));

	QMUX QL_INST_QMUX_BL0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_BL0_padClk));

	QMUX QL_INST_QMUX_BL1 (.GMUXIN(GND),.IS(VCC),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_BL1_tpGCLKBUF));

	QMUX QL_INST_QMUX_BL2 (.GMUXIN(GND),.IS(VCC),.QHSCK(nx22245z2),.IZ(nx22245z2_QMUX_BL2_tpGCLKBUF));

	QMUX QL_INST_QMUX_BR0 (.GMUXIN(CLK_int_0__GMUX_0_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_0__QMUX_BR0_padClk));

	QMUX QL_INST_QMUX_BR1 (.GMUXIN(CLK_int_1__GMUX_1_padClk),.IS(GND),.QHSCK(GND),.IZ(CLK_int_1__QMUX_BR1_padClk));

	QMUX QL_INST_QMUX_BR2 (.GMUXIN(GND),.IS(VCC),.QHSCK(not_RESET_0),.IZ(not_RESET_0_QMUX_BR2_tpGCLKBUF));

	QPMUX QL_INST_QMUX_BR3 (.GMUXIN(GND),.IS0(VCC),.IS1(VCC),.QCLKIN(GND),.QHSCK(nx3850z2),.IZ(nx3850z2_QMUX_BR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSTL0_padClk));

	SQEMUX QL_INST_SQMUX_TLSTL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TL1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx34006z2),.IZ(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTL3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx42928z2),.IZ(nx42928z2_SQMUX_TLSTL3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTL4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx39840z1),.IZ(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTL5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(p0_fsm[0]),.IZ(p0_fsm_0__SQMUX_TLSTL5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSTR0_padClk));

	SQEMUX QL_INST_SQMUX_TLSTR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TL1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSTR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx15998z1),.IZ(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTR3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(tcdm_valid_p0_int),.IZ(tcdm_valid_p0_int_SQMUX_TLSTR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSTR4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx32231z2),.IZ(nx32231z2_SQMUX_TLSTR4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSBL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSBL0_padClk));

	SQEMUX QL_INST_SQMUX_TLSBL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TL1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TLSBL1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSBL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx44608z1),.IZ(nx44608z1_SQMUX_TLSBL2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBL3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_73),.IZ(NET_73_SQMUX_TLSBL3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBL4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(lint_ADDR_int[11]),.IZ(lint_ADDR_int_11__SQMUX_TLSBL4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBL5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_75),.IZ(NET_75_SQMUX_TLSBL5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSBR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TL0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TLSBR0_padClk));

	SQEMUX QL_INST_SQMUX_TLSBR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TL1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TLSBR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_33),.IZ(NET_33_SQMUX_TLSBR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBR3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_126),.IZ(NET_126_SQMUX_TLSBR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBR4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_127),.IZ(NET_127_SQMUX_TLSBR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TLSBR5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_30),.IZ(NET_30_SQMUX_TLSBR5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSTL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSTL0_padClk));

	SQEMUX QL_INST_SQMUX_TRSTL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSTL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx11313z1),.IZ(nx11313z1_SQMUX_TRSTL2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTL3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx41193z2),.IZ(nx41193z2_SQMUX_TRSTL3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTL4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(p1_fsm[0]),.IZ(p1_fsm_0__SQMUX_TRSTL4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTL5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_59),.IZ(NET_59_SQMUX_TRSTL5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSTR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSTR0_padClk));

	SQEMUX QL_INST_SQMUX_TRSTR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSTR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx25587z2),.IZ(nx25587z2_SQMUX_TRSTR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTR3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx11312z1),.IZ(nx11312z1_SQMUX_TRSTR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTR4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx36058z2),.IZ(nx36058z2_SQMUX_TRSTR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSTR5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx39177z2),.IZ(nx39177z2_SQMUX_TRSTR5_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBL0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSBL0_padClk));

	SQEMUX QL_INST_SQMUX_TRSBL1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBL2 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_2__QMUX_TR2_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_2__SQMUX_TRSBL2_padClk));

	SQMUX QL_INST_SQMUX_TRSBL3 (.QMUXIN(CLK_int_3__QMUX_TR3_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_3__SQMUX_TRSBL3_padClk));

	SQMUX QL_INST_SQMUX_TRSBL4 (.QMUXIN(CLK_int_4__QMUX_TR4_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_4__SQMUX_TRSBL4_padClk));

	SQMUX QL_INST_SQMUX_TRSBL5 (.QMUXIN(CLK_int_5__QMUX_TR5_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_5__SQMUX_TRSBL5_padClk));

	SQEMUX QL_INST_SQMUX_TRSBR0 (.DEN(GND),.DYNEN(GND),.QMUXIN(CLK_int_0__QMUX_TR0_padClk),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_TRSBR0_padClk));

	SQEMUX QL_INST_SQMUX_TRSBR1 (.DEN(GND),.DYNEN(GND),.QMUXIN(not_RESET_0_QMUX_TR1_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_TRSBR2 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx13970z2),.IZ(nx13970z2_SQMUX_TRSBR2_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBR3 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx12973z2),.IZ(nx12973z2_SQMUX_TRSBR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBR4 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx11312z1),.IZ(nx11312z1_SQMUX_TRSBR4_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_TRSBR5 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx36058z2),.IZ(nx36058z2_SQMUX_TRSBR5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTL0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSTL0_padClk));

	SQMUX QL_INST_SQMUX_BLSTL1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTL2 (.QMUXIN(nx22245z2_QMUX_BL2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(nx22245z2_SQMUX_BLSTL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTL3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx4939z1),.IZ(nx4939z1_SQMUX_BLSTL3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTL4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx12783z2),.IZ(nx12783z2_SQMUX_BLSTL4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTL5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx9707z1),.IZ(nx9707z1_SQMUX_BLSTL5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTR0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSTR0_padClk));

	SQMUX QL_INST_SQMUX_BLSTR1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSTR2 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(tcdm_valid_p2_int),.IZ(tcdm_valid_p2_int_SQMUX_BLSTR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(lint_ADDR_int[2]),.IZ(lint_ADDR_int_2__SQMUX_BLSTR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_21),.IZ(NET_21_SQMUX_BLSTR4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSTR5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_27),.IZ(NET_27_SQMUX_BLSTR5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBL0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSBL0_padClk));

	SQMUX QL_INST_SQMUX_BLSBL1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBL2 (.QMUXIN(nx22245z2_QMUX_BL2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(nx22245z2_SQMUX_BLSBL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBL3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_482),.IZ(NET_482_SQMUX_BLSBL3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBL4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(p2_fsm[0]),.IZ(p2_fsm_0__SQMUX_BLSBL4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBL5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(p2_fsm[4]),.IZ(p2_fsm_4__SQMUX_BLSBL5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBR0 (.QMUXIN(CLK_int_0__QMUX_BL0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BLSBR0_padClk));

	SQMUX QL_INST_SQMUX_BLSBR1 (.QMUXIN(not_RESET_0_QMUX_BL1_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BLSBR2 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx33579z1),.IZ(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BLSBR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx14650z1),.IZ(nx14650z1_SQMUX_BLSBR3_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTL0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSTL0_padClk));

	SQMUX QL_INST_SQMUX_BRSTL1 (.QMUXIN(CLK_int_1__QMUX_BR1_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_1__SQMUX_BRSTL1_padClk));

	SQMUX QL_INST_SQMUX_BRSTL2 (.QMUXIN(not_RESET_0_QMUX_BR2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSTL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTL3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_62),.IZ(NET_62_SQMUX_BRSTL3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTL4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(apb_fsm[0]),.IZ(apb_fsm_0__SQMUX_BRSTL4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTL5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(lint_ADDR_int[13]),.IZ(lint_ADDR_int_13__SQMUX_BRSTL5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTR0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSTR0_padClk));

	SQMUX QL_INST_SQMUX_BRSTR1 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(nx63842z2),.IZ(nx63842z2_SQMUX_BRSTR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSTR2 (.QMUXIN(not_RESET_0_QMUX_BR2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSTR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx40548z2),.IZ(nx40548z2_SQMUX_BRSTR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx60851z2),.IZ(nx60851z2_SQMUX_BRSTR4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSTR5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx60936z2),.IZ(nx60936z2_SQMUX_BRSTR5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSBL0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSBL0_padClk));

	SQMUX QL_INST_SQMUX_BRSBL1 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(p3_fsm[0]),.IZ(p3_fsm_0__SQMUX_BRSBL1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSBL2 (.QMUXIN(not_RESET_0_QMUX_BR2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSBL2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBL3 (.DEN(GND),.DYNEN(GND),.QMUXIN(nx3850z2_QMUX_BR3_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(nx3850z2_SQMUX_BRSBL3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBL4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(NET_113),.IZ(NET_113_SQMUX_BRSBL4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBL5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx11311z1),.IZ(nx11311z1_SQMUX_BRSBL5_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSBR0 (.QMUXIN(CLK_int_0__QMUX_BR0_padClk),.SELECT(GND),.SQHSCK(GND),.IZ(CLK_int_0__SQMUX_BRSBR0_padClk));

	SQMUX QL_INST_SQMUX_BRSBR1 (.QMUXIN(GND),.SELECT(VCC),.SQHSCK(NET_0),.IZ(NET_0_SQMUX_BRSBR1_tpGCLKBUF));

	SQMUX QL_INST_SQMUX_BRSBR2 (.QMUXIN(not_RESET_0_QMUX_BR2_tpGCLKBUF),.SELECT(GND),.SQHSCK(GND),.IZ(not_RESET_0_SQMUX_BRSBR2_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBR3 (.DEN(GND),.DYNEN(GND),.QMUXIN(nx3850z2_QMUX_BR3_tpGCLKBUF),.SELECT(GND),.SEN(VCC),.SQHSCK(GND),.IZ(nx3850z2_SQMUX_BRSBR3_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBR4 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx25788z3),.IZ(nx25788z3_SQMUX_BRSBR4_tpGCLKBUF));

	SQEMUX QL_INST_SQMUX_BRSBR5 (.DEN(GND),.DYNEN(GND),.QMUXIN(GND),.SELECT(VCC),.SEN(VCC),.SQHSCK(nx3786z2),.IZ(nx3786z2_SQMUX_BRSBR5_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSTL_1 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_1_padClk));

	CAND QL_INST_CAND0_TLSTL_2 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_2_padClk));

	CAND QL_INST_CAND0_TLSTL_3 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_3_padClk));

	CAND QL_INST_CAND0_TLSTL_4 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_4_padClk));

	CAND QL_INST_CAND0_TLSTL_5 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_5_padClk));

	CAND QL_INST_CAND0_TLSTL_6 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_6_padClk));

	CAND QL_INST_CAND0_TLSTL_7 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_7_padClk));

	CAND QL_INST_CAND0_TLSTL_8 (.CLKIN(CLK_int_0__SQMUX_TLSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTL_8_padClk));

	CAND QL_INST_CAND1_TLSTL_1 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_1_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_2 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_2_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_3 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_3_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_4 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_4_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_5 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_6 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_6_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_7 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_7_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTL_8 (.CLKIN(not_RESET_0_SQMUX_TLSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTL_8_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_4 (.CLKIN(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z2_CAND2_TLSTL_4_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_5 (.CLKIN(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z2_CAND2_TLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_6 (.CLKIN(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z2_CAND2_TLSTL_6_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_7 (.CLKIN(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z2_CAND2_TLSTL_7_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTL_8 (.CLKIN(nx34006z2_SQMUX_TLSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx34006z2_CAND2_TLSTL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_4 (.CLKIN(nx42928z2_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx42928z2_CAND3_TLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_5 (.CLKIN(nx42928z2_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx42928z2_CAND3_TLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_6 (.CLKIN(nx42928z2_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx42928z2_CAND3_TLSTL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_7 (.CLKIN(nx42928z2_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx42928z2_CAND3_TLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTL_8 (.CLKIN(nx42928z2_SQMUX_TLSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx42928z2_CAND3_TLSTL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_1 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_2 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_3 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTL_4 (.CLKIN(nx39840z1_SQMUX_TLSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39840z1_CAND4_TLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTL_7 (.CLKIN(p0_fsm_0__SQMUX_TLSTL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(p0_fsm_0__CAND5_TLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSTL_8 (.CLKIN(p0_fsm_0__SQMUX_TLSTL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(p0_fsm_0__CAND5_TLSTL_8_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSTR_9 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_9_padClk));

	CAND QL_INST_CAND0_TLSTR_10 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_10_padClk));

	CAND QL_INST_CAND0_TLSTR_11 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_11_padClk));

	CAND QL_INST_CAND0_TLSTR_12 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_12_padClk));

	CAND QL_INST_CAND0_TLSTR_13 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_13_padClk));

	CAND QL_INST_CAND0_TLSTR_14 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_14_padClk));

	CAND QL_INST_CAND0_TLSTR_15 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_15_padClk));

	CAND QL_INST_CAND0_TLSTR_16 (.CLKIN(CLK_int_0__SQMUX_TLSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSTR_16_padClk));

	CAND QL_INST_CAND1_TLSTR_9 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_9_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_10 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_10_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_11 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_12 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_13 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_14 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_15 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_15_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSTR_16 (.CLKIN(not_RESET_0_SQMUX_TLSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSTR_16_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_11 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_12 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_13 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSTR_14 (.CLKIN(nx15998z1_SQMUX_TLSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx15998z1_CAND2_TLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_9 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND3_TLSTR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_10 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND3_TLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_13 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND3_TLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_14 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND3_TLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_15 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND3_TLSTR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSTR_16 (.CLKIN(tcdm_valid_p0_int_SQMUX_TLSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p0_int_CAND3_TLSTR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_14 (.CLKIN(nx32231z2_SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx32231z2_CAND4_TLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSTR_15 (.CLKIN(nx32231z2_SQMUX_TLSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx32231z2_CAND4_TLSTR_15_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSBL_0 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_0_padClk));

	CAND QL_INST_CAND0_TLSBL_1 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_1_padClk));

	CAND QL_INST_CAND0_TLSBL_2 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_2_padClk));

	CAND QL_INST_CAND0_TLSBL_3 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_3_padClk));

	CAND QL_INST_CAND0_TLSBL_4 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_4_padClk));

	CAND QL_INST_CAND0_TLSBL_5 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_5_padClk));

	CAND QL_INST_CAND0_TLSBL_6 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_6_padClk));

	CAND QL_INST_CAND0_TLSBL_7 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_7_padClk));

	CAND QL_INST_CAND0_TLSBL_8 (.CLKIN(CLK_int_0__SQMUX_TLSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBL_8_padClk));

	CAND QL_INST_CAND1_TLSBL_1 (.CLKIN(not_RESET_0_SQMUX_TLSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBL_1_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBL_2 (.CLKIN(not_RESET_0_SQMUX_TLSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBL_2_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBL_3 (.CLKIN(not_RESET_0_SQMUX_TLSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBL_3_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBL_4 (.CLKIN(not_RESET_0_SQMUX_TLSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBL_4_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBL_5 (.CLKIN(not_RESET_0_SQMUX_TLSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBL_5_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBL_6 (.CLKIN(not_RESET_0_SQMUX_TLSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBL_6_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBL_7 (.CLKIN(not_RESET_0_SQMUX_TLSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBL_7_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBL_8 (.CLKIN(not_RESET_0_SQMUX_TLSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBL_8_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_1 (.CLKIN(nx44608z1_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(nx44608z1_CAND2_TLSBL_1_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_2 (.CLKIN(nx44608z1_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(nx44608z1_CAND2_TLSBL_2_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_3 (.CLKIN(nx44608z1_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(nx44608z1_CAND2_TLSBL_3_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_4 (.CLKIN(nx44608z1_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(nx44608z1_CAND2_TLSBL_4_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBL_5 (.CLKIN(nx44608z1_SQMUX_TLSBL2_tpGCLKBUF),.SEN(VCC),.IZ(nx44608z1_CAND2_TLSBL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_1 (.CLKIN(NET_73_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_73_CAND3_TLSBL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_2 (.CLKIN(NET_73_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_73_CAND3_TLSBL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_3 (.CLKIN(NET_73_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_73_CAND3_TLSBL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBL_4 (.CLKIN(NET_73_SQMUX_TLSBL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_73_CAND3_TLSBL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBL_1 (.CLKIN(lint_ADDR_int_11__SQMUX_TLSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_11__CAND4_TLSBL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBL_2 (.CLKIN(lint_ADDR_int_11__SQMUX_TLSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_11__CAND4_TLSBL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBL_6 (.CLKIN(lint_ADDR_int_11__SQMUX_TLSBL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(lint_ADDR_int_11__CAND4_TLSBL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBL_1 (.CLKIN(NET_75_SQMUX_TLSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_75_CAND5_TLSBL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBL_2 (.CLKIN(NET_75_SQMUX_TLSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_75_CAND5_TLSBL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBL_3 (.CLKIN(NET_75_SQMUX_TLSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_75_CAND5_TLSBL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBL_6 (.CLKIN(NET_75_SQMUX_TLSBL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_75_CAND5_TLSBL_6_tpGCLKBUF));

	CAND QL_INST_CAND0_TLSBR_9 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_9_padClk));

	CAND QL_INST_CAND0_TLSBR_10 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_10_padClk));

	CAND QL_INST_CAND0_TLSBR_11 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_11_padClk));

	CAND QL_INST_CAND0_TLSBR_12 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_12_padClk));

	CAND QL_INST_CAND0_TLSBR_13 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_13_padClk));

	CAND QL_INST_CAND0_TLSBR_14 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_14_padClk));

	CAND QL_INST_CAND0_TLSBR_15 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_15_padClk));

	CAND QL_INST_CAND0_TLSBR_16 (.CLKIN(CLK_int_0__SQMUX_TLSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TLSBR_16_padClk));

	CAND QL_INST_CAND1_TLSBR_9 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_9_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_10 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_10_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_11 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_11_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_12 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_12_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_13 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_13_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_14 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_15 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_15_tpGCLKBUF));

	CAND QL_INST_CAND1_TLSBR_16 (.CLKIN(not_RESET_0_SQMUX_TLSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TLSBR_16_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_10 (.CLKIN(NET_33_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(NET_33_CAND2_TLSBR_10_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_11 (.CLKIN(NET_33_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(NET_33_CAND2_TLSBR_11_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_12 (.CLKIN(NET_33_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(NET_33_CAND2_TLSBR_12_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_14 (.CLKIN(NET_33_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(NET_33_CAND2_TLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND2_TLSBR_16 (.CLKIN(NET_33_SQMUX_TLSBR2_tpGCLKBUF),.SEN(VCC),.IZ(NET_33_CAND2_TLSBR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_10 (.CLKIN(NET_126_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_126_CAND3_TLSBR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_11 (.CLKIN(NET_126_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_126_CAND3_TLSBR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_12 (.CLKIN(NET_126_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_126_CAND3_TLSBR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_13 (.CLKIN(NET_126_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_126_CAND3_TLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TLSBR_14 (.CLKIN(NET_126_SQMUX_TLSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_126_CAND3_TLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_9 (.CLKIN(NET_127_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_127_CAND4_TLSBR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_10 (.CLKIN(NET_127_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_127_CAND4_TLSBR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_12 (.CLKIN(NET_127_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_127_CAND4_TLSBR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_13 (.CLKIN(NET_127_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_127_CAND4_TLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_14 (.CLKIN(NET_127_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_127_CAND4_TLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TLSBR_15 (.CLKIN(NET_127_SQMUX_TLSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_127_CAND4_TLSBR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBR_10 (.CLKIN(NET_30_SQMUX_TLSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_30_CAND5_TLSBR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TLSBR_11 (.CLKIN(NET_30_SQMUX_TLSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_30_CAND5_TLSBR_11_tpGCLKBUF));

	CAND QL_INST_CAND0_TRSTL_17 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_17_padClk));

	CAND QL_INST_CAND0_TRSTL_18 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_18_padClk));

	CAND QL_INST_CAND0_TRSTL_19 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_19_padClk));

	CAND QL_INST_CAND0_TRSTL_20 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_20_padClk));

	CAND QL_INST_CAND0_TRSTL_21 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_21_padClk));

	CAND QL_INST_CAND0_TRSTL_22 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_22_padClk));

	CAND QL_INST_CAND0_TRSTL_23 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_23_padClk));

	CAND QL_INST_CAND0_TRSTL_24 (.CLKIN(CLK_int_0__SQMUX_TRSTL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTL_24_padClk));

	CAND QL_INST_CAND1_TRSTL_17 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_17_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTL_18 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_18_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTL_19 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_19_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTL_20 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_20_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTL_21 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_21_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTL_22 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_22_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTL_23 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_23_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTL_24 (.CLKIN(not_RESET_0_SQMUX_TRSTL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTL_24_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTL_17 (.CLKIN(nx11313z1_SQMUX_TRSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx11313z1_CAND2_TRSTL_17_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTL_18 (.CLKIN(nx11313z1_SQMUX_TRSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx11313z1_CAND2_TRSTL_18_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTL_19 (.CLKIN(nx11313z1_SQMUX_TRSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx11313z1_CAND2_TRSTL_19_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTL_20 (.CLKIN(nx11313z1_SQMUX_TRSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx11313z1_CAND2_TRSTL_20_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTL_21 (.CLKIN(nx11313z1_SQMUX_TRSTL2_tpGCLKBUF),.SEN(VCC),.IZ(nx11313z1_CAND2_TRSTL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTL_17 (.CLKIN(nx41193z2_SQMUX_TRSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z2_CAND3_TRSTL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTL_18 (.CLKIN(nx41193z2_SQMUX_TRSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z2_CAND3_TRSTL_18_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTL_19 (.CLKIN(nx41193z2_SQMUX_TRSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z2_CAND3_TRSTL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTL_20 (.CLKIN(nx41193z2_SQMUX_TRSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z2_CAND3_TRSTL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTL_21 (.CLKIN(nx41193z2_SQMUX_TRSTL3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx41193z2_CAND3_TRSTL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTL_22 (.CLKIN(p1_fsm_0__SQMUX_TRSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(p1_fsm_0__CAND4_TRSTL_22_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTL_23 (.CLKIN(p1_fsm_0__SQMUX_TRSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(p1_fsm_0__CAND4_TRSTL_23_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTL_24 (.CLKIN(p1_fsm_0__SQMUX_TRSTL4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(p1_fsm_0__CAND4_TRSTL_24_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSTL_19 (.CLKIN(NET_59_SQMUX_TRSTL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_59_CAND5_TRSTL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSTL_20 (.CLKIN(NET_59_SQMUX_TRSTL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_59_CAND5_TRSTL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSTL_21 (.CLKIN(NET_59_SQMUX_TRSTL5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_59_CAND5_TRSTL_21_tpGCLKBUF));

	CAND QL_INST_CAND0_TRSTR_25 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_25_padClk));

	CAND QL_INST_CAND0_TRSTR_26 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_26_padClk));

	CAND QL_INST_CAND0_TRSTR_27 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_27_padClk));

	CAND QL_INST_CAND0_TRSTR_28 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_28_padClk));

	CAND QL_INST_CAND0_TRSTR_29 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_29_padClk));

	CAND QL_INST_CAND0_TRSTR_33 (.CLKIN(CLK_int_0__SQMUX_TRSTR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSTR_33_padClk));

	CAND QL_INST_CAND1_TRSTR_25 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_25_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_26 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_26_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_27 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_27_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_28 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_28_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSTR_29 (.CLKIN(not_RESET_0_SQMUX_TRSTR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSTR_29_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTR_25 (.CLKIN(nx25587z2_SQMUX_TRSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx25587z2_CAND2_TRSTR_25_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSTR_26 (.CLKIN(nx25587z2_SQMUX_TRSTR2_tpGCLKBUF),.SEN(VCC),.IZ(nx25587z2_CAND2_TRSTR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_25 (.CLKIN(nx11312z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx11312z1_CAND3_TRSTR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_26 (.CLKIN(nx11312z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx11312z1_CAND3_TRSTR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_27 (.CLKIN(nx11312z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx11312z1_CAND3_TRSTR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_28 (.CLKIN(nx11312z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx11312z1_CAND3_TRSTR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSTR_29 (.CLKIN(nx11312z1_SQMUX_TRSTR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx11312z1_CAND3_TRSTR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_25 (.CLKIN(nx36058z2_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx36058z2_CAND4_TRSTR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_26 (.CLKIN(nx36058z2_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx36058z2_CAND4_TRSTR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_27 (.CLKIN(nx36058z2_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx36058z2_CAND4_TRSTR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_28 (.CLKIN(nx36058z2_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx36058z2_CAND4_TRSTR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSTR_29 (.CLKIN(nx36058z2_SQMUX_TRSTR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx36058z2_CAND4_TRSTR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSTR_25 (.CLKIN(nx39177z2_SQMUX_TRSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39177z2_CAND5_TRSTR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSTR_26 (.CLKIN(nx39177z2_SQMUX_TRSTR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx39177z2_CAND5_TRSTR_26_tpGCLKBUF));

	CAND QL_INST_CAND0_TRSBL_17 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_17_padClk));

	CAND QL_INST_CAND0_TRSBL_18 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_18_padClk));

	CAND QL_INST_CAND0_TRSBL_19 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_19_padClk));

	CAND QL_INST_CAND0_TRSBL_21 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_21_padClk));

	CAND QL_INST_CAND0_TRSBL_22 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_22_padClk));

	CAND QL_INST_CAND0_TRSBL_23 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_23_padClk));

	CAND QL_INST_CAND0_TRSBL_24 (.CLKIN(CLK_int_0__SQMUX_TRSBL0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBL_24_padClk));

	CAND QL_INST_CAND1_TRSBL_17 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_17_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_18 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_18_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_19 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_19_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_21 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_21_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_22 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_22_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_23 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_23_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBL_24 (.CLKIN(not_RESET_0_SQMUX_TRSBL1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBL_24_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBL_18 (.CLKIN(CLK_int_2__SQMUX_TRSBL2_padClk),.SEN(VCC),.IZ(CLK_int_2__CAND2_TRSBL_18_padClk));

	CANDEN QL_INST_CAND3_TRSBL_17 (.CLKIN(CLK_int_3__SQMUX_TRSBL3_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_3__CAND3_TRSBL_17_padClk));

	CANDEN QL_INST_CAND4_TRSBL_20 (.CLKIN(CLK_int_4__SQMUX_TRSBL4_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_4__CAND4_TRSBL_20_padClk));

	CANDEN QL_INST_CAND5_TRSBL_17 (.CLKIN(CLK_int_5__SQMUX_TRSBL5_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_5__CAND5_TRSBL_17_padClk));

	CAND QL_INST_CAND0_TRSBR_25 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_25_padClk));

	CAND QL_INST_CAND0_TRSBR_26 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_26_padClk));

	CAND QL_INST_CAND0_TRSBR_27 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_27_padClk));

	CAND QL_INST_CAND0_TRSBR_28 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_28_padClk));

	CAND QL_INST_CAND0_TRSBR_29 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_29_padClk));

	CAND QL_INST_CAND0_TRSBR_33 (.CLKIN(CLK_int_0__SQMUX_TRSBR0_padClk),.SEN(VCC),.IZ(CLK_int_0__CAND0_TRSBR_33_padClk));

	CAND QL_INST_CAND1_TRSBR_25 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_25_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBR_26 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_26_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBR_27 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_27_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBR_28 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_28_tpGCLKBUF));

	CAND QL_INST_CAND1_TRSBR_29 (.CLKIN(not_RESET_0_SQMUX_TRSBR1_tpGCLKBUF),.SEN(VCC),.IZ(not_RESET_0_CAND1_TRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_26 (.CLKIN(nx13970z2_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx13970z2_CAND2_TRSBR_26_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_27 (.CLKIN(nx13970z2_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx13970z2_CAND2_TRSBR_27_tpGCLKBUF));

	CAND QL_INST_CAND2_TRSBR_28 (.CLKIN(nx13970z2_SQMUX_TRSBR2_tpGCLKBUF),.SEN(VCC),.IZ(nx13970z2_CAND2_TRSBR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBR_26 (.CLKIN(nx12973z2_SQMUX_TRSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx12973z2_CAND3_TRSBR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND3_TRSBR_27 (.CLKIN(nx12973z2_SQMUX_TRSBR3_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx12973z2_CAND3_TRSBR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBR_25 (.CLKIN(nx11312z1_SQMUX_TRSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx11312z1_CAND4_TRSBR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBR_26 (.CLKIN(nx11312z1_SQMUX_TRSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx11312z1_CAND4_TRSBR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBR_27 (.CLKIN(nx11312z1_SQMUX_TRSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx11312z1_CAND4_TRSBR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBR_28 (.CLKIN(nx11312z1_SQMUX_TRSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx11312z1_CAND4_TRSBR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND4_TRSBR_29 (.CLKIN(nx11312z1_SQMUX_TRSBR4_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx11312z1_CAND4_TRSBR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBR_25 (.CLKIN(nx36058z2_SQMUX_TRSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx36058z2_CAND5_TRSBR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBR_26 (.CLKIN(nx36058z2_SQMUX_TRSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx36058z2_CAND5_TRSBR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBR_27 (.CLKIN(nx36058z2_SQMUX_TRSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx36058z2_CAND5_TRSBR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBR_28 (.CLKIN(nx36058z2_SQMUX_TRSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx36058z2_CAND5_TRSBR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND5_TRSBR_29 (.CLKIN(nx36058z2_SQMUX_TRSBR5_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx36058z2_CAND5_TRSBR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSTL_1 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_1_padClk));

	CANDEN QL_INST_CAND0_BLSTL_2 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_2_padClk));

	CANDEN QL_INST_CAND0_BLSTL_3 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_3_padClk));

	CANDEN QL_INST_CAND0_BLSTL_4 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_4_padClk));

	CANDEN QL_INST_CAND0_BLSTL_5 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_5_padClk));

	CANDEN QL_INST_CAND0_BLSTL_6 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_6_padClk));

	CANDEN QL_INST_CAND0_BLSTL_7 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_7_padClk));

	CANDEN QL_INST_CAND0_BLSTL_8 (.CLKIN(CLK_int_0__SQMUX_BLSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTL_8_padClk));

	CANDEN QL_INST_CAND1_BLSTL_1 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_2 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_3 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_3_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_4 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_4_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_5 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_6 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_7 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTL_8 (.CLKIN(not_RESET_0_SQMUX_BLSTL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_5 (.CLKIN(nx22245z2_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx22245z2_CAND2_BLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_6 (.CLKIN(nx22245z2_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx22245z2_CAND2_BLSTL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_7 (.CLKIN(nx22245z2_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx22245z2_CAND2_BLSTL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTL_8 (.CLKIN(nx22245z2_SQMUX_BLSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx22245z2_CAND2_BLSTL_8_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTL_1 (.CLKIN(nx4939z1_SQMUX_BLSTL3_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND3_BLSTL_1_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTL_2 (.CLKIN(nx4939z1_SQMUX_BLSTL3_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND3_BLSTL_2_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTL_3 (.CLKIN(nx4939z1_SQMUX_BLSTL3_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND3_BLSTL_3_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTL_4 (.CLKIN(nx4939z1_SQMUX_BLSTL3_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND3_BLSTL_4_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTL_5 (.CLKIN(nx4939z1_SQMUX_BLSTL3_tpGCLKBUF),.SEN(VCC),.IZ(nx4939z1_CAND3_BLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTL_5 (.CLKIN(nx12783z2_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(nx12783z2_CAND4_BLSTL_5_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTL_6 (.CLKIN(nx12783z2_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(nx12783z2_CAND4_BLSTL_6_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTL_7 (.CLKIN(nx12783z2_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(nx12783z2_CAND4_BLSTL_7_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTL_8 (.CLKIN(nx12783z2_SQMUX_BLSTL4_tpGCLKBUF),.SEN(VCC),.IZ(nx12783z2_CAND4_BLSTL_8_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_1 (.CLKIN(nx9707z1_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(nx9707z1_CAND5_BLSTL_1_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_2 (.CLKIN(nx9707z1_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(nx9707z1_CAND5_BLSTL_2_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_3 (.CLKIN(nx9707z1_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(nx9707z1_CAND5_BLSTL_3_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTL_5 (.CLKIN(nx9707z1_SQMUX_BLSTL5_tpGCLKBUF),.SEN(VCC),.IZ(nx9707z1_CAND5_BLSTL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSTR_9 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_9_padClk));

	CANDEN QL_INST_CAND0_BLSTR_10 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_10_padClk));

	CANDEN QL_INST_CAND0_BLSTR_11 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_11_padClk));

	CANDEN QL_INST_CAND0_BLSTR_12 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_12_padClk));

	CANDEN QL_INST_CAND0_BLSTR_13 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_13_padClk));

	CANDEN QL_INST_CAND0_BLSTR_14 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_14_padClk));

	CANDEN QL_INST_CAND0_BLSTR_15 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_15_padClk));

	CANDEN QL_INST_CAND0_BLSTR_16 (.CLKIN(CLK_int_0__SQMUX_BLSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSTR_16_padClk));

	CANDEN QL_INST_CAND1_BLSTR_9 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_10 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_11 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_12 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_13 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_14 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_15 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSTR_16 (.CLKIN(not_RESET_0_SQMUX_BLSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSTR_16_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_10 (.CLKIN(tcdm_valid_p2_int_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p2_int_CAND2_BLSTR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_12 (.CLKIN(tcdm_valid_p2_int_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p2_int_CAND2_BLSTR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_13 (.CLKIN(tcdm_valid_p2_int_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p2_int_CAND2_BLSTR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSTR_15 (.CLKIN(tcdm_valid_p2_int_SQMUX_BLSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(tcdm_valid_p2_int_CAND2_BLSTR_15_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_11 (.CLKIN(lint_ADDR_int_2__SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(lint_ADDR_int_2__CAND3_BLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_12 (.CLKIN(lint_ADDR_int_2__SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(lint_ADDR_int_2__CAND3_BLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_14 (.CLKIN(lint_ADDR_int_2__SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(lint_ADDR_int_2__CAND3_BLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_15 (.CLKIN(lint_ADDR_int_2__SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(lint_ADDR_int_2__CAND3_BLSTR_15_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSTR_16 (.CLKIN(lint_ADDR_int_2__SQMUX_BLSTR3_tpGCLKBUF),.SEN(VCC),.IZ(lint_ADDR_int_2__CAND3_BLSTR_16_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_12 (.CLKIN(NET_21_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_21_CAND4_BLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_13 (.CLKIN(NET_21_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_21_CAND4_BLSTR_13_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSTR_15 (.CLKIN(NET_21_SQMUX_BLSTR4_tpGCLKBUF),.SEN(VCC),.IZ(NET_21_CAND4_BLSTR_15_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_10 (.CLKIN(NET_27_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_27_CAND5_BLSTR_10_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_11 (.CLKIN(NET_27_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_27_CAND5_BLSTR_11_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_12 (.CLKIN(NET_27_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_27_CAND5_BLSTR_12_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_14 (.CLKIN(NET_27_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_27_CAND5_BLSTR_14_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSTR_15 (.CLKIN(NET_27_SQMUX_BLSTR5_tpGCLKBUF),.SEN(VCC),.IZ(NET_27_CAND5_BLSTR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSBL_1 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_1_padClk));

	CANDEN QL_INST_CAND0_BLSBL_2 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_2_padClk));

	CANDEN QL_INST_CAND0_BLSBL_5 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_5_padClk));

	CANDEN QL_INST_CAND0_BLSBL_6 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_6_padClk));

	CANDEN QL_INST_CAND0_BLSBL_7 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_7_padClk));

	CANDEN QL_INST_CAND0_BLSBL_8 (.CLKIN(CLK_int_0__SQMUX_BLSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBL_8_padClk));

	CANDEN QL_INST_CAND1_BLSBL_1 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_1_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_2 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_2_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_5 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_6 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_7 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBL_8 (.CLKIN(not_RESET_0_SQMUX_BLSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_5 (.CLKIN(nx22245z2_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx22245z2_CAND2_BLSBL_5_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_6 (.CLKIN(nx22245z2_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx22245z2_CAND2_BLSBL_6_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_7 (.CLKIN(nx22245z2_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx22245z2_CAND2_BLSBL_7_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBL_8 (.CLKIN(nx22245z2_SQMUX_BLSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx22245z2_CAND2_BLSBL_8_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBL_5 (.CLKIN(NET_482_SQMUX_BLSBL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_482_CAND3_BLSBL_5_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBL_6 (.CLKIN(NET_482_SQMUX_BLSBL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_482_CAND3_BLSBL_6_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBL_8 (.CLKIN(NET_482_SQMUX_BLSBL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_482_CAND3_BLSBL_8_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBL_6 (.CLKIN(p2_fsm_0__SQMUX_BLSBL4_tpGCLKBUF),.SEN(VCC),.IZ(p2_fsm_0__CAND4_BLSBL_6_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBL_7 (.CLKIN(p2_fsm_0__SQMUX_BLSBL4_tpGCLKBUF),.SEN(VCC),.IZ(p2_fsm_0__CAND4_BLSBL_7_tpGCLKBUF));

	CAND QL_INST_CAND4_BLSBL_8 (.CLKIN(p2_fsm_0__SQMUX_BLSBL4_tpGCLKBUF),.SEN(VCC),.IZ(p2_fsm_0__CAND4_BLSBL_8_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSBL_5 (.CLKIN(p2_fsm_4__SQMUX_BLSBL5_tpGCLKBUF),.SEN(VCC),.IZ(p2_fsm_4__CAND5_BLSBL_5_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSBL_6 (.CLKIN(p2_fsm_4__SQMUX_BLSBL5_tpGCLKBUF),.SEN(VCC),.IZ(p2_fsm_4__CAND5_BLSBL_6_tpGCLKBUF));

	CAND QL_INST_CAND5_BLSBL_8 (.CLKIN(p2_fsm_4__SQMUX_BLSBL5_tpGCLKBUF),.SEN(VCC),.IZ(p2_fsm_4__CAND5_BLSBL_8_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BLSBR_9 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_9_padClk));

	CANDEN QL_INST_CAND0_BLSBR_10 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_10_padClk));

	CANDEN QL_INST_CAND0_BLSBR_11 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_11_padClk));

	CANDEN QL_INST_CAND0_BLSBR_12 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_12_padClk));

	CANDEN QL_INST_CAND0_BLSBR_13 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_13_padClk));

	CANDEN QL_INST_CAND0_BLSBR_14 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_14_padClk));

	CANDEN QL_INST_CAND0_BLSBR_15 (.CLKIN(CLK_int_0__SQMUX_BLSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BLSBR_15_padClk));

	CANDEN QL_INST_CAND1_BLSBR_9 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_9_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_10 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_10_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_11 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_12 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_13 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_14 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_14_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BLSBR_15 (.CLKIN(not_RESET_0_SQMUX_BLSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND1_BLSBR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_11 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_11_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_12 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_12_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_13 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_13_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BLSBR_14 (.CLKIN(nx33579z1_SQMUX_BLSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx33579z1_CAND2_BLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_14 (.CLKIN(nx14650z1_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx14650z1_CAND3_BLSBR_14_tpGCLKBUF));

	CAND QL_INST_CAND3_BLSBR_15 (.CLKIN(nx14650z1_SQMUX_BLSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx14650z1_CAND3_BLSBR_15_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSTL_17 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_17_padClk));

	CANDEN QL_INST_CAND0_BRSTL_18 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_18_padClk));

	CANDEN QL_INST_CAND0_BRSTL_19 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_19_padClk));

	CANDEN QL_INST_CAND0_BRSTL_20 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_20_padClk));

	CANDEN QL_INST_CAND0_BRSTL_21 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_21_padClk));

	CANDEN QL_INST_CAND0_BRSTL_22 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_22_padClk));

	CANDEN QL_INST_CAND0_BRSTL_23 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_23_padClk));

	CANDEN QL_INST_CAND0_BRSTL_24 (.CLKIN(CLK_int_0__SQMUX_BRSTL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTL_24_padClk));

	CANDEN QL_INST_CAND1_BRSTL_20 (.CLKIN(CLK_int_1__SQMUX_BRSTL1_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_1__CAND1_BRSTL_20_padClk));

	CANDEN QL_INST_CAND1_BRSTL_21 (.CLKIN(CLK_int_1__SQMUX_BRSTL1_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_1__CAND1_BRSTL_21_padClk));

	CANDEN QL_INST_CAND2_BRSTL_17 (.CLKIN(not_RESET_0_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_18 (.CLKIN(not_RESET_0_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTL_18_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_19 (.CLKIN(not_RESET_0_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_20 (.CLKIN(not_RESET_0_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_21 (.CLKIN(not_RESET_0_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_22 (.CLKIN(not_RESET_0_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTL_22_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_23 (.CLKIN(not_RESET_0_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTL_23_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTL_24 (.CLKIN(not_RESET_0_SQMUX_BRSTL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTL_24_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTL_17 (.CLKIN(NET_62_SQMUX_BRSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_62_CAND3_BRSTL_17_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTL_18 (.CLKIN(NET_62_SQMUX_BRSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_62_CAND3_BRSTL_18_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTL_19 (.CLKIN(NET_62_SQMUX_BRSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_62_CAND3_BRSTL_19_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTL_20 (.CLKIN(NET_62_SQMUX_BRSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_62_CAND3_BRSTL_20_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTL_21 (.CLKIN(NET_62_SQMUX_BRSTL3_tpGCLKBUF),.SEN(VCC),.IZ(NET_62_CAND3_BRSTL_21_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTL_17 (.CLKIN(apb_fsm_0__SQMUX_BRSTL4_tpGCLKBUF),.SEN(VCC),.IZ(apb_fsm_0__CAND4_BRSTL_17_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTL_18 (.CLKIN(apb_fsm_0__SQMUX_BRSTL4_tpGCLKBUF),.SEN(VCC),.IZ(apb_fsm_0__CAND4_BRSTL_18_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTL_19 (.CLKIN(apb_fsm_0__SQMUX_BRSTL4_tpGCLKBUF),.SEN(VCC),.IZ(apb_fsm_0__CAND4_BRSTL_19_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTL_20 (.CLKIN(apb_fsm_0__SQMUX_BRSTL4_tpGCLKBUF),.SEN(VCC),.IZ(apb_fsm_0__CAND4_BRSTL_20_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSTL_18 (.CLKIN(lint_ADDR_int_13__SQMUX_BRSTL5_tpGCLKBUF),.SEN(VCC),.IZ(lint_ADDR_int_13__CAND5_BRSTL_18_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSTL_19 (.CLKIN(lint_ADDR_int_13__SQMUX_BRSTL5_tpGCLKBUF),.SEN(VCC),.IZ(lint_ADDR_int_13__CAND5_BRSTL_19_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSTL_20 (.CLKIN(lint_ADDR_int_13__SQMUX_BRSTL5_tpGCLKBUF),.SEN(VCC),.IZ(lint_ADDR_int_13__CAND5_BRSTL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSTR_25 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_25_padClk));

	CANDEN QL_INST_CAND0_BRSTR_26 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_26_padClk));

	CANDEN QL_INST_CAND0_BRSTR_27 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_27_padClk));

	CANDEN QL_INST_CAND0_BRSTR_28 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_28_padClk));

	CANDEN QL_INST_CAND0_BRSTR_29 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_29_padClk));

	CANDEN QL_INST_CAND0_BRSTR_33 (.CLKIN(CLK_int_0__SQMUX_BRSTR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSTR_33_padClk));

	CANDEN QL_INST_CAND1_BRSTR_25 (.CLKIN(nx63842z2_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx63842z2_CAND1_BRSTR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTR_26 (.CLKIN(nx63842z2_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx63842z2_CAND1_BRSTR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTR_27 (.CLKIN(nx63842z2_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx63842z2_CAND1_BRSTR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSTR_28 (.CLKIN(nx63842z2_SQMUX_BRSTR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(nx63842z2_CAND1_BRSTR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_25 (.CLKIN(not_RESET_0_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_26 (.CLKIN(not_RESET_0_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_27 (.CLKIN(not_RESET_0_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_28 (.CLKIN(not_RESET_0_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSTR_29 (.CLKIN(not_RESET_0_SQMUX_BRSTR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSTR_29_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTR_25 (.CLKIN(nx40548z2_SQMUX_BRSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx40548z2_CAND3_BRSTR_25_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTR_26 (.CLKIN(nx40548z2_SQMUX_BRSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx40548z2_CAND3_BRSTR_26_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSTR_27 (.CLKIN(nx40548z2_SQMUX_BRSTR3_tpGCLKBUF),.SEN(VCC),.IZ(nx40548z2_CAND3_BRSTR_27_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTR_27 (.CLKIN(nx60851z2_SQMUX_BRSTR4_tpGCLKBUF),.SEN(VCC),.IZ(nx60851z2_CAND4_BRSTR_27_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSTR_28 (.CLKIN(nx60851z2_SQMUX_BRSTR4_tpGCLKBUF),.SEN(VCC),.IZ(nx60851z2_CAND4_BRSTR_28_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSTR_25 (.CLKIN(nx60936z2_SQMUX_BRSTR5_tpGCLKBUF),.SEN(VCC),.IZ(nx60936z2_CAND5_BRSTR_25_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSTR_26 (.CLKIN(nx60936z2_SQMUX_BRSTR5_tpGCLKBUF),.SEN(VCC),.IZ(nx60936z2_CAND5_BRSTR_26_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSTR_27 (.CLKIN(nx60936z2_SQMUX_BRSTR5_tpGCLKBUF),.SEN(VCC),.IZ(nx60936z2_CAND5_BRSTR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSBL_17 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_17_padClk));

	CANDEN QL_INST_CAND0_BRSBL_18 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_18_padClk));

	CANDEN QL_INST_CAND0_BRSBL_19 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_19_padClk));

	CANDEN QL_INST_CAND0_BRSBL_20 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_20_padClk));

	CANDEN QL_INST_CAND0_BRSBL_21 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_21_padClk));

	CANDEN QL_INST_CAND0_BRSBL_22 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_22_padClk));

	CANDEN QL_INST_CAND0_BRSBL_23 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_23_padClk));

	CANDEN QL_INST_CAND0_BRSBL_24 (.CLKIN(CLK_int_0__SQMUX_BRSBL0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBL_24_padClk));

	CANDEN QL_INST_CAND1_BRSBL_21 (.CLKIN(p3_fsm_0__SQMUX_BRSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(p3_fsm_0__CAND1_BRSBL_21_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBL_22 (.CLKIN(p3_fsm_0__SQMUX_BRSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(p3_fsm_0__CAND1_BRSBL_22_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBL_23 (.CLKIN(p3_fsm_0__SQMUX_BRSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(p3_fsm_0__CAND1_BRSBL_23_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBL_24 (.CLKIN(p3_fsm_0__SQMUX_BRSBL1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(p3_fsm_0__CAND1_BRSBL_24_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBL_17 (.CLKIN(not_RESET_0_SQMUX_BRSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBL_17_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBL_18 (.CLKIN(not_RESET_0_SQMUX_BRSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBL_18_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBL_19 (.CLKIN(not_RESET_0_SQMUX_BRSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBL_19_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBL_20 (.CLKIN(not_RESET_0_SQMUX_BRSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBL_23 (.CLKIN(not_RESET_0_SQMUX_BRSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBL_23_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBL_24 (.CLKIN(not_RESET_0_SQMUX_BRSBL2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBL_24_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBL_23 (.CLKIN(nx3850z2_SQMUX_BRSBL3_tpGCLKBUF),.SEN(VCC),.IZ(nx3850z2_CAND3_BRSBL_23_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBL_24 (.CLKIN(nx3850z2_SQMUX_BRSBL3_tpGCLKBUF),.SEN(VCC),.IZ(nx3850z2_CAND3_BRSBL_24_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBL_17 (.CLKIN(NET_113_SQMUX_BRSBL4_tpGCLKBUF),.SEN(VCC),.IZ(NET_113_CAND4_BRSBL_17_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBL_18 (.CLKIN(NET_113_SQMUX_BRSBL4_tpGCLKBUF),.SEN(VCC),.IZ(NET_113_CAND4_BRSBL_18_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBL_19 (.CLKIN(NET_113_SQMUX_BRSBL4_tpGCLKBUF),.SEN(VCC),.IZ(NET_113_CAND4_BRSBL_19_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBL_20 (.CLKIN(NET_113_SQMUX_BRSBL4_tpGCLKBUF),.SEN(VCC),.IZ(NET_113_CAND4_BRSBL_20_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBL_17 (.CLKIN(nx11311z1_SQMUX_BRSBL5_tpGCLKBUF),.SEN(VCC),.IZ(nx11311z1_CAND5_BRSBL_17_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBL_18 (.CLKIN(nx11311z1_SQMUX_BRSBL5_tpGCLKBUF),.SEN(VCC),.IZ(nx11311z1_CAND5_BRSBL_18_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBL_19 (.CLKIN(nx11311z1_SQMUX_BRSBL5_tpGCLKBUF),.SEN(VCC),.IZ(nx11311z1_CAND5_BRSBL_19_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBL_20 (.CLKIN(nx11311z1_SQMUX_BRSBL5_tpGCLKBUF),.SEN(VCC),.IZ(nx11311z1_CAND5_BRSBL_20_tpGCLKBUF));

	CANDEN QL_INST_CAND0_BRSBR_25 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_25_padClk));

	CANDEN QL_INST_CAND0_BRSBR_26 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_26_padClk));

	CANDEN QL_INST_CAND0_BRSBR_27 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_27_padClk));

	CANDEN QL_INST_CAND0_BRSBR_28 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_28_padClk));

	CANDEN QL_INST_CAND0_BRSBR_29 (.CLKIN(CLK_int_0__SQMUX_BRSBR0_padClk),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(CLK_int_0__CAND0_BRSBR_29_padClk));

	CANDEN QL_INST_CAND1_BRSBR_25 (.CLKIN(NET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_0_CAND1_BRSBR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_26 (.CLKIN(NET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_0_CAND1_BRSBR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_27 (.CLKIN(NET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_0_CAND1_BRSBR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_28 (.CLKIN(NET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_0_CAND1_BRSBR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND1_BRSBR_29 (.CLKIN(NET_0_SQMUX_BRSBR1_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(NET_0_CAND1_BRSBR_29_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_25 (.CLKIN(not_RESET_0_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBR_25_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_26 (.CLKIN(not_RESET_0_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBR_26_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_27 (.CLKIN(not_RESET_0_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBR_27_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_28 (.CLKIN(not_RESET_0_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBR_28_tpGCLKBUF));

	CANDEN QL_INST_CAND2_BRSBR_29 (.CLKIN(not_RESET_0_SQMUX_BRSBR2_tpGCLKBUF),.DEN(GND),.DYNEN(GND),.SEN(VCC),.IZ(not_RESET_0_CAND2_BRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_25 (.CLKIN(nx3850z2_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx3850z2_CAND3_BRSBR_25_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_26 (.CLKIN(nx3850z2_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx3850z2_CAND3_BRSBR_26_tpGCLKBUF));

	CAND QL_INST_CAND3_BRSBR_27 (.CLKIN(nx3850z2_SQMUX_BRSBR3_tpGCLKBUF),.SEN(VCC),.IZ(nx3850z2_CAND3_BRSBR_27_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBR_25 (.CLKIN(nx25788z3_SQMUX_BRSBR4_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z3_CAND4_BRSBR_25_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBR_26 (.CLKIN(nx25788z3_SQMUX_BRSBR4_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z3_CAND4_BRSBR_26_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBR_27 (.CLKIN(nx25788z3_SQMUX_BRSBR4_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z3_CAND4_BRSBR_27_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBR_28 (.CLKIN(nx25788z3_SQMUX_BRSBR4_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z3_CAND4_BRSBR_28_tpGCLKBUF));

	CAND QL_INST_CAND4_BRSBR_29 (.CLKIN(nx25788z3_SQMUX_BRSBR4_tpGCLKBUF),.SEN(VCC),.IZ(nx25788z3_CAND4_BRSBR_29_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBR_25 (.CLKIN(nx3786z2_SQMUX_BRSBR5_tpGCLKBUF),.SEN(VCC),.IZ(nx3786z2_CAND5_BRSBR_25_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBR_26 (.CLKIN(nx3786z2_SQMUX_BRSBR5_tpGCLKBUF),.SEN(VCC),.IZ(nx3786z2_CAND5_BRSBR_26_tpGCLKBUF));

	CAND QL_INST_CAND5_BRSBR_27 (.CLKIN(nx3786z2_SQMUX_BRSBR5_tpGCLKBUF),.SEN(VCC),.IZ(nx3786z2_CAND5_BRSBR_27_tpGCLKBUF));

	qlOBUF QL_INST_F2A_T_1_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTL_1_padClk),.OUT_OBUF(m1_oper0_rclk));

	qlOBUF QL_INST_F2A_T_1_1 (.IN_OBUF(CLK_int_0__CAND0_TLSTL_1_padClk),.OUT_OBUF(m1_oper1_rclk));

	qlOBUF QL_INST_F2A_T_1_4 (.IN_OBUF(CLK_int_0__CAND0_TLSTL_1_padClk),.OUT_OBUF(m0_coef_wclk));

	qlOBUF QL_INST_F2A_T_2_0 (.IN_OBUF(CLK_int_0__CAND0_TLSTL_2_padClk),.OUT_OBUF(m0_oper0_rclk));

	qlOBUF QL_INST_F2A_T_2_1 (.IN_OBUF(m0_oper0_wmode_dup_0[1]),.OUT_OBUF(m0_oper0_wmode[1]));

	qlOBUF QL_INST_F2A_T_2_2 (.IN_OBUF(m0_oper0_wmode_dup_0[0]),.OUT_OBUF(m0_oper0_wmode[0]));

	qlOBUF QL_INST_F2A_T_2_4 (.IN_OBUF(m0_oper0_rmode_dup_0[1]),.OUT_OBUF(m0_oper0_rmode[1]));

	qlOBUF QL_INST_F2A_T_2_5 (.IN_OBUF(m0_oper0_rmode_dup_0[0]),.OUT_OBUF(m0_oper0_rmode[0]));

	qlOBUF QL_INST_F2A_T_2_6 (.IN_OBUF(m0_oper0_wdata_dup_0[31]),.OUT_OBUF(m0_oper0_wdata[31]));

	qlOBUF QL_INST_F2A_T_2_7 (.IN_OBUF(m0_oper0_wdata_dup_0[30]),.OUT_OBUF(m0_oper0_wdata[30]));

	qlOBUF QL_INST_F2A_T_2_8 (.IN_OBUF(m0_oper0_wdata_dup_0[29]),.OUT_OBUF(m0_oper0_wdata[29]));

	qlOBUF QL_INST_F2A_T_2_9 (.IN_OBUF(m0_oper0_wdata_dup_0[28]),.OUT_OBUF(m0_oper0_wdata[28]));

	qlOBUF QL_INST_F2A_T_2_10 (.IN_OBUF(m0_oper0_wdata_dup_0[27]),.OUT_OBUF(m0_oper0_wdata[27]));

	qlOBUF QL_INST_F2A_T_2_11 (.IN_OBUF(m0_oper0_wdata_dup_0[26]),.OUT_OBUF(m0_oper0_wdata[26]));

	qlOBUF QL_INST_F2A_T_2_12 (.IN_OBUF(m0_oper0_wdata_dup_0[25]),.OUT_OBUF(m0_oper0_wdata[25]));

	qlOBUF QL_INST_F2A_T_2_13 (.IN_OBUF(m0_oper0_wdata_dup_0[24]),.OUT_OBUF(m0_oper0_wdata[24]));

	qlOBUF QL_INST_F2A_T_2_14 (.IN_OBUF(m0_oper0_wdata_dup_0[23]),.OUT_OBUF(m0_oper0_wdata[23]));

	qlOBUF QL_INST_F2A_T_2_15 (.IN_OBUF(m0_oper0_wdata_dup_0[22]),.OUT_OBUF(m0_oper0_wdata[22]));

	qlOBUF QL_INST_F2A_T_2_16 (.IN_OBUF(m0_oper0_wdata_dup_0[21]),.OUT_OBUF(m0_oper0_wdata[21]));

	qlOBUF QL_INST_F2A_T_2_17 (.IN_OBUF(m0_oper0_wdata_dup_0[20]),.OUT_OBUF(m0_oper0_wdata[20]));

	qlIBUF QL_INST_A2F_T_2_0 (.IN_IBUF(m0_oper0_rdata[31]),.OUT_IBUF(m0_oper0_rdata_int[31]));

	qlIBUF QL_INST_A2F_T_2_1 (.IN_IBUF(m0_oper0_rdata[30]),.OUT_IBUF(m0_oper0_rdata_int[30]));

	qlIBUF QL_INST_A2F_T_2_2 (.IN_IBUF(m0_oper0_rdata[29]),.OUT_IBUF(m0_oper0_rdata_int[29]));

	qlIBUF QL_INST_A2F_T_2_3 (.IN_IBUF(m0_oper0_rdata[28]),.OUT_IBUF(m0_oper0_rdata_int[28]));

	qlOBUF QL_INST_F2A_T_3_0 (.IN_OBUF(m0_oper0_wdata_dup_0[19]),.OUT_OBUF(m0_oper0_wdata[19]));

	qlOBUF QL_INST_F2A_T_3_1 (.IN_OBUF(m0_oper0_wdata_dup_0[18]),.OUT_OBUF(m0_oper0_wdata[18]));

	qlOBUF QL_INST_F2A_T_3_2 (.IN_OBUF(m0_oper0_wdata_dup_0[17]),.OUT_OBUF(m0_oper0_wdata[17]));

	qlOBUF QL_INST_F2A_T_3_3 (.IN_OBUF(m0_oper0_wdata_dup_0[16]),.OUT_OBUF(m0_oper0_wdata[16]));

	qlOBUF QL_INST_F2A_T_3_4 (.IN_OBUF(m0_oper0_wdata_dup_0[15]),.OUT_OBUF(m0_oper0_wdata[15]));

	qlOBUF QL_INST_F2A_T_3_5 (.IN_OBUF(m0_oper0_wdata_dup_0[14]),.OUT_OBUF(m0_oper0_wdata[14]));

	qlOBUF QL_INST_F2A_T_3_6 (.IN_OBUF(m0_oper0_wdata_dup_0[13]),.OUT_OBUF(m0_oper0_wdata[13]));

	qlOBUF QL_INST_F2A_T_3_7 (.IN_OBUF(m0_oper0_wdata_dup_0[12]),.OUT_OBUF(m0_oper0_wdata[12]));

	qlOBUF QL_INST_F2A_T_3_8 (.IN_OBUF(m0_oper0_wdata_dup_0[11]),.OUT_OBUF(m0_oper0_wdata[11]));

	qlOBUF QL_INST_F2A_T_3_9 (.IN_OBUF(m0_oper0_wdata_dup_0[10]),.OUT_OBUF(m0_oper0_wdata[10]));

	qlOBUF QL_INST_F2A_T_3_10 (.IN_OBUF(m0_oper0_wdata_dup_0[9]),.OUT_OBUF(m0_oper0_wdata[9]));

	qlOBUF QL_INST_F2A_T_3_11 (.IN_OBUF(m0_oper0_wdata_dup_0[8]),.OUT_OBUF(m0_oper0_wdata[8]));

	qlIBUF QL_INST_A2F_T_3_0 (.IN_IBUF(m0_oper0_rdata[27]),.OUT_IBUF(m0_oper0_rdata_int[27]));

	qlIBUF QL_INST_A2F_T_3_1 (.IN_IBUF(m0_oper0_rdata[26]),.OUT_IBUF(m0_oper0_rdata_int[26]));

	qlIBUF QL_INST_A2F_T_3_2 (.IN_IBUF(m0_oper0_rdata[25]),.OUT_IBUF(m0_oper0_rdata_int[25]));

	qlIBUF QL_INST_A2F_T_3_3 (.IN_IBUF(m0_oper0_rdata[24]),.OUT_IBUF(m0_oper0_rdata_int[24]));

	qlIBUF QL_INST_A2F_T_3_4 (.IN_IBUF(m0_oper0_rdata[23]),.OUT_IBUF(m0_oper0_rdata_int[23]));

	qlIBUF QL_INST_A2F_T_3_5 (.IN_IBUF(m0_oper0_rdata[22]),.OUT_IBUF(m0_oper0_rdata_int[22]));

	qlOBUF QL_INST_F2A_T_4_0 (.IN_OBUF(m0_oper0_wdata_dup_0[7]),.OUT_OBUF(m0_oper0_wdata[7]));

	qlOBUF QL_INST_F2A_T_4_1 (.IN_OBUF(m0_oper0_wdata_dup_0[6]),.OUT_OBUF(m0_oper0_wdata[6]));

	qlOBUF QL_INST_F2A_T_4_2 (.IN_OBUF(m0_oper0_wdata_dup_0[5]),.OUT_OBUF(m0_oper0_wdata[5]));

	qlOBUF QL_INST_F2A_T_4_3 (.IN_OBUF(m0_oper0_wdata_dup_0[4]),.OUT_OBUF(m0_oper0_wdata[4]));

	qlOBUF QL_INST_F2A_T_4_4 (.IN_OBUF(m0_oper0_wdata_dup_0[3]),.OUT_OBUF(m0_oper0_wdata[3]));

	qlOBUF QL_INST_F2A_T_4_5 (.IN_OBUF(m0_oper0_wdata_dup_0[2]),.OUT_OBUF(m0_oper0_wdata[2]));

	qlOBUF QL_INST_F2A_T_4_6 (.IN_OBUF(m0_oper0_wdata_dup_0[1]),.OUT_OBUF(m0_oper0_wdata[1]));

	qlOBUF QL_INST_F2A_T_4_7 (.IN_OBUF(m0_oper0_wdata_dup_0[0]),.OUT_OBUF(m0_oper0_wdata[0]));

	qlOBUF QL_INST_F2A_T_4_8 (.IN_OBUF(m0_oper0_waddr_dup_0[11]),.OUT_OBUF(m0_oper0_waddr[11]));

	qlOBUF QL_INST_F2A_T_4_9 (.IN_OBUF(m0_oper0_waddr_dup_0[10]),.OUT_OBUF(m0_oper0_waddr[10]));

	qlOBUF QL_INST_F2A_T_4_10 (.IN_OBUF(m0_oper0_waddr_dup_0[9]),.OUT_OBUF(m0_oper0_waddr[9]));

	qlOBUF QL_INST_F2A_T_4_11 (.IN_OBUF(m0_oper0_waddr_dup_0[8]),.OUT_OBUF(m0_oper0_waddr[8]));

	qlOBUF QL_INST_F2A_T_4_12 (.IN_OBUF(m0_oper0_waddr_dup_0[7]),.OUT_OBUF(m0_oper0_waddr[7]));

	qlOBUF QL_INST_F2A_T_4_13 (.IN_OBUF(m0_oper0_waddr_dup_0[6]),.OUT_OBUF(m0_oper0_waddr[6]));

	qlOBUF QL_INST_F2A_T_4_14 (.IN_OBUF(m0_oper0_waddr_dup_0[5]),.OUT_OBUF(m0_oper0_waddr[5]));

	qlOBUF QL_INST_F2A_T_4_15 (.IN_OBUF(m0_oper0_waddr_dup_0[4]),.OUT_OBUF(m0_oper0_waddr[4]));

	qlOBUF QL_INST_F2A_T_4_16 (.IN_OBUF(m0_oper0_waddr_dup_0[3]),.OUT_OBUF(m0_oper0_waddr[3]));

	qlOBUF QL_INST_F2A_T_4_17 (.IN_OBUF(m0_oper0_waddr_dup_0[2]),.OUT_OBUF(m0_oper0_waddr[2]));

	qlIBUF QL_INST_A2F_T_4_0 (.IN_IBUF(m0_oper0_rdata[21]),.OUT_IBUF(m0_oper0_rdata_int[21]));

	qlIBUF QL_INST_A2F_T_4_1 (.IN_IBUF(m0_oper0_rdata[20]),.OUT_IBUF(m0_oper0_rdata_int[20]));

	qlIBUF QL_INST_A2F_T_4_2 (.IN_IBUF(m0_oper0_rdata[19]),.OUT_IBUF(m0_oper0_rdata_int[19]));

	qlIBUF QL_INST_A2F_T_4_3 (.IN_IBUF(m0_oper0_rdata[18]),.OUT_IBUF(m0_oper0_rdata_int[18]));

	qlIBUF QL_INST_A2F_T_4_4 (.IN_IBUF(m0_oper0_rdata[17]),.OUT_IBUF(m0_oper0_rdata_int[17]));

	qlIBUF QL_INST_A2F_T_4_5 (.IN_IBUF(m0_oper0_rdata[16]),.OUT_IBUF(m0_oper0_rdata_int[16]));

	qlIBUF QL_INST_A2F_T_4_6 (.IN_IBUF(m0_oper0_rdata[15]),.OUT_IBUF(m0_oper0_rdata_int[15]));

	qlIBUF QL_INST_A2F_T_4_7 (.IN_IBUF(m0_oper0_rdata[14]),.OUT_IBUF(m0_oper0_rdata_int[14]));

	qlOBUF QL_INST_F2A_T_5_0 (.IN_OBUF(m0_oper0_waddr_dup_0[1]),.OUT_OBUF(m0_oper0_waddr[1]));

	qlOBUF QL_INST_F2A_T_5_1 (.IN_OBUF(m0_oper0_waddr_dup_0[0]),.OUT_OBUF(m0_oper0_waddr[0]));

	qlOBUF QL_INST_F2A_T_5_3 (.IN_OBUF(m0_oper0_raddr_dup_0[11]),.OUT_OBUF(m0_oper0_raddr[11]));

	qlOBUF QL_INST_F2A_T_5_4 (.IN_OBUF(m0_oper0_raddr_dup_0[10]),.OUT_OBUF(m0_oper0_raddr[10]));

	qlOBUF QL_INST_F2A_T_5_5 (.IN_OBUF(m0_oper0_raddr_dup_0[9]),.OUT_OBUF(m0_oper0_raddr[9]));

	qlOBUF QL_INST_F2A_T_5_6 (.IN_OBUF(m0_oper0_raddr_dup_0[8]),.OUT_OBUF(m0_oper0_raddr[8]));

	qlOBUF QL_INST_F2A_T_5_7 (.IN_OBUF(m0_oper0_raddr_dup_0[7]),.OUT_OBUF(m0_oper0_raddr[7]));

	qlOBUF QL_INST_F2A_T_5_8 (.IN_OBUF(m0_oper0_raddr_dup_0[6]),.OUT_OBUF(m0_oper0_raddr[6]));

	qlOBUF QL_INST_F2A_T_5_9 (.IN_OBUF(m0_oper0_raddr_dup_0[5]),.OUT_OBUF(m0_oper0_raddr[5]));

	qlOBUF QL_INST_F2A_T_5_10 (.IN_OBUF(m0_oper0_raddr_dup_0[4]),.OUT_OBUF(m0_oper0_raddr[4]));

	qlOBUF QL_INST_F2A_T_5_11 (.IN_OBUF(m0_oper0_raddr_dup_0[3]),.OUT_OBUF(m0_oper0_raddr[3]));

	qlIBUF QL_INST_A2F_T_5_0 (.IN_IBUF(m0_oper0_rdata[13]),.OUT_IBUF(m0_oper0_rdata_int[13]));

	qlIBUF QL_INST_A2F_T_5_1 (.IN_IBUF(m0_oper0_rdata[12]),.OUT_IBUF(m0_oper0_rdata_int[12]));

	qlIBUF QL_INST_A2F_T_5_2 (.IN_IBUF(m0_oper0_rdata[11]),.OUT_IBUF(m0_oper0_rdata_int[11]));

	qlIBUF QL_INST_A2F_T_5_3 (.IN_IBUF(m0_oper0_rdata[10]),.OUT_IBUF(m0_oper0_rdata_int[10]));

	qlIBUF QL_INST_A2F_T_5_4 (.IN_IBUF(m0_oper0_rdata[9]),.OUT_IBUF(m0_oper0_rdata_int[9]));

	qlIBUF QL_INST_A2F_T_5_5 (.IN_IBUF(m0_oper0_rdata[8]),.OUT_IBUF(m0_oper0_rdata_int[8]));

	qlOBUF QL_INST_F2A_T_6_0 (.IN_OBUF(m0_oper0_we_dup_0),.OUT_OBUF(m0_oper0_we));

	qlOBUF QL_INST_F2A_T_6_1 (.IN_OBUF(m0_oper0_raddr_dup_0[2]),.OUT_OBUF(m0_oper0_raddr[2]));

	qlOBUF QL_INST_F2A_T_6_2 (.IN_OBUF(m0_oper0_raddr_dup_0[1]),.OUT_OBUF(m0_oper0_raddr[1]));

	qlOBUF QL_INST_F2A_T_6_3 (.IN_OBUF(m0_oper0_raddr_dup_0[0]),.OUT_OBUF(m0_oper0_raddr[0]));

	qlOBUF QL_INST_F2A_T_6_4 (.IN_OBUF(m1_m0_clr_dup_0),.OUT_OBUF(m1_m0_clr));

	qlOBUF QL_INST_F2A_T_6_5 (.IN_OBUF(m1_m1_sat_dup_0),.OUT_OBUF(m1_m1_sat));

	qlOBUF QL_INST_F2A_T_6_6 (.IN_OBUF(m0_m0_outsel_dup_0[5]),.OUT_OBUF(m0_m0_outsel[5]));

	qlOBUF QL_INST_F2A_T_6_7 (.IN_OBUF(m0_m0_outsel_dup_0[4]),.OUT_OBUF(m0_m0_outsel[4]));

	qlOBUF QL_INST_F2A_T_6_8 (.IN_OBUF(m0_m0_outsel_dup_0[3]),.OUT_OBUF(m0_m0_outsel[3]));

	qlOBUF QL_INST_F2A_T_6_9 (.IN_OBUF(m0_m0_outsel_dup_0[2]),.OUT_OBUF(m0_m0_outsel[2]));

	qlOBUF QL_INST_F2A_T_6_10 (.IN_OBUF(m0_m0_outsel_dup_0[1]),.OUT_OBUF(m0_m0_outsel[1]));

	qlOBUF QL_INST_F2A_T_6_11 (.IN_OBUF(m0_m0_outsel_dup_0[0]),.OUT_OBUF(m0_m0_outsel[0]));

	qlOBUF QL_INST_F2A_T_6_12 (.IN_OBUF(m1_oper0_wdsel_dup_0),.OUT_OBUF(m1_oper0_wdsel));

	qlOBUF QL_INST_F2A_T_6_13 (.IN_OBUF(m1_oper1_wdsel_dup_0),.OUT_OBUF(m1_oper1_wdsel));

	qlOBUF QL_INST_F2A_T_6_14 (.IN_OBUF(m0_oper1_wdsel_dup_0),.OUT_OBUF(m0_oper1_wdsel));

	qlOBUF QL_INST_F2A_T_6_15 (.IN_OBUF(m0_oper0_rdata_int[31]),.OUT_OBUF(m0_m0_oper_in[31]));

	qlOBUF QL_INST_F2A_T_6_16 (.IN_OBUF(m0_oper0_rdata_int[30]),.OUT_OBUF(m0_m0_oper_in[30]));

	qlOBUF QL_INST_F2A_T_6_17 (.IN_OBUF(m0_oper0_rdata_int[29]),.OUT_OBUF(m0_m0_oper_in[29]));

	DBUF QL_INST_F2Adef_T_6_1 (.IN_DBUF(GND),.OUT_DBUF(m1_oper1_powerdn));

	qlIBUF QL_INST_A2F_T_6_0 (.IN_IBUF(m0_oper0_rdata[7]),.OUT_IBUF(m0_oper0_rdata_int[7]));

	qlIBUF QL_INST_A2F_T_6_1 (.IN_IBUF(m0_oper0_rdata[6]),.OUT_IBUF(m0_oper0_rdata_int[6]));

	qlIBUF QL_INST_A2F_T_6_2 (.IN_IBUF(m0_oper0_rdata[5]),.OUT_IBUF(m0_oper0_rdata_int[5]));

	qlIBUF QL_INST_A2F_T_6_3 (.IN_IBUF(m0_oper0_rdata[4]),.OUT_IBUF(m0_oper0_rdata_int[4]));

	qlIBUF QL_INST_A2F_T_6_4 (.IN_IBUF(m0_oper0_rdata[3]),.OUT_IBUF(m0_oper0_rdata_int[3]));

	qlIBUF QL_INST_A2F_T_6_5 (.IN_IBUF(m0_oper0_rdata[2]),.OUT_IBUF(m0_oper0_rdata_int[2]));

	qlIBUF QL_INST_A2F_T_6_6 (.IN_IBUF(m0_oper0_rdata[1]),.OUT_IBUF(m0_oper0_rdata_int[1]));

	qlIBUF QL_INST_A2F_T_6_7 (.IN_IBUF(m0_oper0_rdata[0]),.OUT_IBUF(m0_oper0_rdata_int[0]));

	qlOBUF QL_INST_F2A_T_7_0 (.IN_OBUF(m1_m0_sat_dup_0),.OUT_OBUF(m1_m0_sat));

	qlOBUF QL_INST_F2A_T_7_1 (.IN_OBUF(m0_oper0_rdata_int[28]),.OUT_OBUF(m0_m0_oper_in[28]));

	qlOBUF QL_INST_F2A_T_7_2 (.IN_OBUF(m0_oper0_rdata_int[27]),.OUT_OBUF(m0_m0_oper_in[27]));

	qlOBUF QL_INST_F2A_T_7_3 (.IN_OBUF(m0_oper0_rdata_int[26]),.OUT_OBUF(m0_m0_oper_in[26]));

	qlOBUF QL_INST_F2A_T_7_4 (.IN_OBUF(m0_oper0_rdata_int[25]),.OUT_OBUF(m0_m0_oper_in[25]));

	qlOBUF QL_INST_F2A_T_7_5 (.IN_OBUF(m0_oper0_rdata_int[24]),.OUT_OBUF(m0_m0_oper_in[24]));

	qlOBUF QL_INST_F2A_T_7_6 (.IN_OBUF(m0_oper0_rdata_int[23]),.OUT_OBUF(m0_m0_oper_in[23]));

	qlOBUF QL_INST_F2A_T_7_7 (.IN_OBUF(m0_oper0_rdata_int[22]),.OUT_OBUF(m0_m0_oper_in[22]));

	qlOBUF QL_INST_F2A_T_7_8 (.IN_OBUF(m0_oper0_rdata_int[21]),.OUT_OBUF(m0_m0_oper_in[21]));

	qlOBUF QL_INST_F2A_T_7_9 (.IN_OBUF(m0_oper0_rdata_int[20]),.OUT_OBUF(m0_m0_oper_in[20]));

	qlOBUF QL_INST_F2A_T_7_10 (.IN_OBUF(m0_oper0_rdata_int[19]),.OUT_OBUF(m0_m0_oper_in[19]));

	qlOBUF QL_INST_F2A_T_7_11 (.IN_OBUF(m0_oper0_rdata_int[18]),.OUT_OBUF(m0_m0_oper_in[18]));

	qlIBUF QL_INST_A2F_T_7_0 (.IN_IBUF(m0_m0_dataout[31]),.OUT_IBUF(m0_m0_dataout_int[31]));

	qlIBUF QL_INST_A2F_T_7_1 (.IN_IBUF(m0_m0_dataout[30]),.OUT_IBUF(m0_m0_dataout_int[30]));

	qlIBUF QL_INST_A2F_T_7_2 (.IN_IBUF(m0_m0_dataout[29]),.OUT_IBUF(m0_m0_dataout_int[29]));

	qlIBUF QL_INST_A2F_T_7_3 (.IN_IBUF(m0_m0_dataout[28]),.OUT_IBUF(m0_m0_dataout_int[28]));

	qlIBUF QL_INST_A2F_T_7_4 (.IN_IBUF(m0_m0_dataout[27]),.OUT_IBUF(m0_m0_dataout_int[27]));

	qlIBUF QL_INST_A2F_T_7_5 (.IN_IBUF(m0_m0_dataout[26]),.OUT_IBUF(m0_m0_dataout_int[26]));

	qlOBUF QL_INST_F2A_T_8_0 (.IN_OBUF(m0_oper0_rdata_int[17]),.OUT_OBUF(m0_m0_oper_in[17]));

	qlOBUF QL_INST_F2A_T_8_1 (.IN_OBUF(m0_oper0_rdata_int[16]),.OUT_OBUF(m0_m0_oper_in[16]));

	qlOBUF QL_INST_F2A_T_8_2 (.IN_OBUF(m0_oper0_rdata_int[15]),.OUT_OBUF(m0_m0_oper_in[15]));

	qlOBUF QL_INST_F2A_T_8_3 (.IN_OBUF(m0_oper0_rdata_int[14]),.OUT_OBUF(m0_m0_oper_in[14]));

	qlOBUF QL_INST_F2A_T_8_4 (.IN_OBUF(m0_oper0_rdata_int[13]),.OUT_OBUF(m0_m0_oper_in[13]));

	qlOBUF QL_INST_F2A_T_8_5 (.IN_OBUF(m0_oper0_rdata_int[12]),.OUT_OBUF(m0_m0_oper_in[12]));

	qlOBUF QL_INST_F2A_T_8_6 (.IN_OBUF(m0_oper0_rdata_int[11]),.OUT_OBUF(m0_m0_oper_in[11]));

	qlOBUF QL_INST_F2A_T_8_7 (.IN_OBUF(m0_oper0_rdata_int[10]),.OUT_OBUF(m0_m0_oper_in[10]));

	qlOBUF QL_INST_F2A_T_8_8 (.IN_OBUF(m0_oper0_rdata_int[9]),.OUT_OBUF(m0_m0_oper_in[9]));

	qlOBUF QL_INST_F2A_T_8_9 (.IN_OBUF(m0_oper0_rdata_int[8]),.OUT_OBUF(m0_m0_oper_in[8]));

	qlOBUF QL_INST_F2A_T_8_10 (.IN_OBUF(m0_oper0_rdata_int[7]),.OUT_OBUF(m0_m0_oper_in[7]));

	qlOBUF QL_INST_F2A_T_8_11 (.IN_OBUF(m0_oper0_rdata_int[6]),.OUT_OBUF(m0_m0_oper_in[6]));

	qlOBUF QL_INST_F2A_T_8_12 (.IN_OBUF(m0_oper0_rdata_int[5]),.OUT_OBUF(m0_m0_oper_in[5]));

	qlOBUF QL_INST_F2A_T_8_13 (.IN_OBUF(m0_oper0_rdata_int[4]),.OUT_OBUF(m0_m0_oper_in[4]));

	qlOBUF QL_INST_F2A_T_8_14 (.IN_OBUF(m0_oper0_rdata_int[3]),.OUT_OBUF(m0_m0_oper_in[3]));

	qlOBUF QL_INST_F2A_T_8_15 (.IN_OBUF(m0_oper0_rdata_int[2]),.OUT_OBUF(m0_m0_oper_in[2]));

	qlOBUF QL_INST_F2A_T_8_16 (.IN_OBUF(m0_oper0_rdata_int[1]),.OUT_OBUF(m0_m0_oper_in[1]));

	qlOBUF QL_INST_F2A_T_8_17 (.IN_OBUF(m0_oper0_rdata_int[0]),.OUT_OBUF(m0_m0_oper_in[0]));

	qlIBUF QL_INST_A2F_T_8_0 (.IN_IBUF(m0_m0_dataout[25]),.OUT_IBUF(m0_m0_dataout_int[25]));

	qlIBUF QL_INST_A2F_T_8_1 (.IN_IBUF(m0_m0_dataout[24]),.OUT_IBUF(m0_m0_dataout_int[24]));

	qlIBUF QL_INST_A2F_T_8_2 (.IN_IBUF(m0_m0_dataout[23]),.OUT_IBUF(m0_m0_dataout_int[23]));

	qlIBUF QL_INST_A2F_T_8_3 (.IN_IBUF(m0_m0_dataout[22]),.OUT_IBUF(m0_m0_dataout_int[22]));

	qlIBUF QL_INST_A2F_T_8_4 (.IN_IBUF(m0_m0_dataout[21]),.OUT_IBUF(m0_m0_dataout_int[21]));

	qlIBUF QL_INST_A2F_T_8_5 (.IN_IBUF(m0_m0_dataout[20]),.OUT_IBUF(m0_m0_dataout_int[20]));

	qlIBUF QL_INST_A2F_T_8_6 (.IN_IBUF(m0_m0_dataout[19]),.OUT_IBUF(m0_m0_dataout_int[19]));

	qlIBUF QL_INST_A2F_T_8_7 (.IN_IBUF(m0_m0_dataout[18]),.OUT_IBUF(m0_m0_dataout_int[18]));

	qlOBUF QL_INST_F2A_T_9_0 (.IN_OBUF(m0_m1_clr_dup_0),.OUT_OBUF(m0_m1_clr));

	qlOBUF QL_INST_F2A_T_9_1 (.IN_OBUF(m0_coef_rdata_int[31]),.OUT_OBUF(m0_m0_coef_in[31]));

	qlOBUF QL_INST_F2A_T_9_2 (.IN_OBUF(m0_coef_rdata_int[30]),.OUT_OBUF(m0_m0_coef_in[30]));

	qlOBUF QL_INST_F2A_T_9_3 (.IN_OBUF(m0_coef_rdata_int[29]),.OUT_OBUF(m0_m0_coef_in[29]));

	qlOBUF QL_INST_F2A_T_9_4 (.IN_OBUF(m0_coef_rdata_int[28]),.OUT_OBUF(m0_m0_coef_in[28]));

	qlOBUF QL_INST_F2A_T_9_5 (.IN_OBUF(m0_coef_rdata_int[27]),.OUT_OBUF(m0_m0_coef_in[27]));

	qlOBUF QL_INST_F2A_T_9_6 (.IN_OBUF(m0_coef_rdata_int[26]),.OUT_OBUF(m0_m0_coef_in[26]));

	qlOBUF QL_INST_F2A_T_9_7 (.IN_OBUF(m0_coef_rdata_int[25]),.OUT_OBUF(m0_m0_coef_in[25]));

	qlOBUF QL_INST_F2A_T_9_8 (.IN_OBUF(m0_coef_rdata_int[24]),.OUT_OBUF(m0_m0_coef_in[24]));

	qlOBUF QL_INST_F2A_T_9_9 (.IN_OBUF(m0_coef_rdata_int[23]),.OUT_OBUF(m0_m0_coef_in[23]));

	qlOBUF QL_INST_F2A_T_9_10 (.IN_OBUF(m0_coef_rdata_int[22]),.OUT_OBUF(m0_m0_coef_in[22]));

	qlOBUF QL_INST_F2A_T_9_11 (.IN_OBUF(m0_coef_rdata_int[21]),.OUT_OBUF(m0_m0_coef_in[21]));

	qlIBUF QL_INST_A2F_T_9_0 (.IN_IBUF(m0_m0_dataout[17]),.OUT_IBUF(m0_m0_dataout_int[17]));

	qlIBUF QL_INST_A2F_T_9_1 (.IN_IBUF(m0_m0_dataout[16]),.OUT_IBUF(m0_m0_dataout_int[16]));

	qlIBUF QL_INST_A2F_T_9_2 (.IN_IBUF(m0_m0_dataout[15]),.OUT_IBUF(m0_m0_dataout_int[15]));

	qlIBUF QL_INST_A2F_T_9_3 (.IN_IBUF(m0_m0_dataout[14]),.OUT_IBUF(m0_m0_dataout_int[14]));

	qlIBUF QL_INST_A2F_T_9_4 (.IN_IBUF(m0_m0_dataout[13]),.OUT_IBUF(m0_m0_dataout_int[13]));

	qlIBUF QL_INST_A2F_T_9_5 (.IN_IBUF(m0_m0_dataout[12]),.OUT_IBUF(m0_m0_dataout_int[12]));

	qlOBUF QL_INST_F2A_T_10_0 (.IN_OBUF(m0_coef_rdata_int[20]),.OUT_OBUF(m0_m0_coef_in[20]));

	qlOBUF QL_INST_F2A_T_10_1 (.IN_OBUF(m0_coef_rdata_int[19]),.OUT_OBUF(m0_m0_coef_in[19]));

	qlOBUF QL_INST_F2A_T_10_2 (.IN_OBUF(m0_coef_rdata_int[18]),.OUT_OBUF(m0_m0_coef_in[18]));

	qlOBUF QL_INST_F2A_T_10_3 (.IN_OBUF(m0_coef_rdata_int[17]),.OUT_OBUF(m0_m0_coef_in[17]));

	qlOBUF QL_INST_F2A_T_10_4 (.IN_OBUF(m0_coef_rdata_int[16]),.OUT_OBUF(m0_m0_coef_in[16]));

	qlOBUF QL_INST_F2A_T_10_5 (.IN_OBUF(m0_coef_rdata_int[15]),.OUT_OBUF(m0_m0_coef_in[15]));

	qlOBUF QL_INST_F2A_T_10_6 (.IN_OBUF(m0_coef_rdata_int[14]),.OUT_OBUF(m0_m0_coef_in[14]));

	qlOBUF QL_INST_F2A_T_10_7 (.IN_OBUF(m0_coef_rdata_int[13]),.OUT_OBUF(m0_m0_coef_in[13]));

	qlOBUF QL_INST_F2A_T_10_8 (.IN_OBUF(m0_coef_rdata_int[12]),.OUT_OBUF(m0_m0_coef_in[12]));

	qlOBUF QL_INST_F2A_T_10_9 (.IN_OBUF(m0_coef_rdata_int[11]),.OUT_OBUF(m0_m0_coef_in[11]));

	qlOBUF QL_INST_F2A_T_10_10 (.IN_OBUF(m0_coef_rdata_int[10]),.OUT_OBUF(m0_m0_coef_in[10]));

	qlOBUF QL_INST_F2A_T_10_11 (.IN_OBUF(m0_coef_rdata_int[9]),.OUT_OBUF(m0_m0_coef_in[9]));

	qlOBUF QL_INST_F2A_T_10_12 (.IN_OBUF(m0_coef_rdata_int[8]),.OUT_OBUF(m0_m0_coef_in[8]));

	qlOBUF QL_INST_F2A_T_10_13 (.IN_OBUF(m0_coef_rdata_int[7]),.OUT_OBUF(m0_m0_coef_in[7]));

	qlOBUF QL_INST_F2A_T_10_14 (.IN_OBUF(m0_coef_rdata_int[6]),.OUT_OBUF(m0_m0_coef_in[6]));

	qlOBUF QL_INST_F2A_T_10_15 (.IN_OBUF(m0_coef_rdata_int[5]),.OUT_OBUF(m0_m0_coef_in[5]));

	qlOBUF QL_INST_F2A_T_10_16 (.IN_OBUF(m0_coef_rdata_int[4]),.OUT_OBUF(m0_m0_coef_in[4]));

	qlOBUF QL_INST_F2A_T_10_17 (.IN_OBUF(m0_coef_rdata_int[3]),.OUT_OBUF(m0_m0_coef_in[3]));

	qlIBUF QL_INST_A2F_T_10_0 (.IN_IBUF(m0_m0_dataout[11]),.OUT_IBUF(m0_m0_dataout_int[11]));

	qlIBUF QL_INST_A2F_T_10_1 (.IN_IBUF(m0_m0_dataout[10]),.OUT_IBUF(m0_m0_dataout_int[10]));

	qlIBUF QL_INST_A2F_T_10_2 (.IN_IBUF(m0_m0_dataout[9]),.OUT_IBUF(m0_m0_dataout_int[9]));

	qlIBUF QL_INST_A2F_T_10_3 (.IN_IBUF(m0_m0_dataout[8]),.OUT_IBUF(m0_m0_dataout_int[8]));

	qlIBUF QL_INST_A2F_T_10_4 (.IN_IBUF(m0_m0_dataout[7]),.OUT_IBUF(m0_m0_dataout_int[7]));

	qlIBUF QL_INST_A2F_T_10_5 (.IN_IBUF(m0_m0_dataout[6]),.OUT_IBUF(m0_m0_dataout_int[6]));

	qlIBUF QL_INST_A2F_T_10_6 (.IN_IBUF(m0_m0_dataout[5]),.OUT_IBUF(m0_m0_dataout_int[5]));

	qlIBUF QL_INST_A2F_T_10_7 (.IN_IBUF(m0_m0_dataout[4]),.OUT_IBUF(m0_m0_dataout_int[4]));

	qlOBUF QL_INST_F2A_T_11_0 (.IN_OBUF(m0_coef_rdata_int[2]),.OUT_OBUF(m0_m0_coef_in[2]));

	qlOBUF QL_INST_F2A_T_11_1 (.IN_OBUF(m0_coef_rdata_int[1]),.OUT_OBUF(m0_m0_coef_in[1]));

	qlOBUF QL_INST_F2A_T_11_2 (.IN_OBUF(m0_coef_rdata_int[0]),.OUT_OBUF(m0_m0_coef_in[0]));

	qlOBUF QL_INST_F2A_T_11_3 (.IN_OBUF(m0_m0_mode_dup_0[1]),.OUT_OBUF(m0_m0_mode[1]));

	qlOBUF QL_INST_F2A_T_11_4 (.IN_OBUF(m0_m0_mode_dup_0[0]),.OUT_OBUF(m0_m0_mode[0]));

	qlOBUF QL_INST_F2A_T_11_5 (.IN_OBUF(m0_m1_tc_dup_0),.OUT_OBUF(m0_m1_tc));

	qlOBUF QL_INST_F2A_T_11_6 (.IN_OBUF(m1_m1_reset_dup_0),.OUT_OBUF(m1_m1_reset));

	qlOBUF QL_INST_F2A_T_11_7 (.IN_OBUF(m0_coef_wdata_dup_0[31]),.OUT_OBUF(m0_coef_wdata[31]));

	qlOBUF QL_INST_F2A_T_11_8 (.IN_OBUF(m0_coef_wdata_dup_0[30]),.OUT_OBUF(m0_coef_wdata[30]));

	qlOBUF QL_INST_F2A_T_11_9 (.IN_OBUF(m0_coef_wdata_dup_0[29]),.OUT_OBUF(m0_coef_wdata[29]));

	qlOBUF QL_INST_F2A_T_11_10 (.IN_OBUF(m0_coef_wdata_dup_0[28]),.OUT_OBUF(m0_coef_wdata[28]));

	qlOBUF QL_INST_F2A_T_11_11 (.IN_OBUF(m0_coef_wdata_dup_0[27]),.OUT_OBUF(m0_coef_wdata[27]));

	qlIBUF QL_INST_A2F_T_11_0 (.IN_IBUF(m0_m0_dataout[3]),.OUT_IBUF(m0_m0_dataout_int[3]));

	qlIBUF QL_INST_A2F_T_11_1 (.IN_IBUF(m0_m0_dataout[2]),.OUT_IBUF(m0_m0_dataout_int[2]));

	qlIBUF QL_INST_A2F_T_11_2 (.IN_IBUF(m0_m0_dataout[1]),.OUT_IBUF(m0_m0_dataout_int[1]));

	qlIBUF QL_INST_A2F_T_11_3 (.IN_IBUF(m0_m0_dataout[0]),.OUT_IBUF(m0_m0_dataout_int[0]));

	qlIBUF QL_INST_A2F_T_11_4 (.IN_IBUF(m0_coef_rdata[31]),.OUT_IBUF(m0_coef_rdata_int[31]));

	qlIBUF QL_INST_A2F_T_11_5 (.IN_IBUF(m0_coef_rdata[30]),.OUT_IBUF(m0_coef_rdata_int[30]));

	qlOBUF QL_INST_F2A_T_12_0 (.IN_OBUF(m0_coef_wdata_dup_0[26]),.OUT_OBUF(m0_coef_wdata[26]));

	qlOBUF QL_INST_F2A_T_12_1 (.IN_OBUF(m0_coef_wdata_dup_0[25]),.OUT_OBUF(m0_coef_wdata[25]));

	qlOBUF QL_INST_F2A_T_12_2 (.IN_OBUF(m0_coef_wdata_dup_0[24]),.OUT_OBUF(m0_coef_wdata[24]));

	qlOBUF QL_INST_F2A_T_12_3 (.IN_OBUF(m0_coef_wdata_dup_0[23]),.OUT_OBUF(m0_coef_wdata[23]));

	qlOBUF QL_INST_F2A_T_12_4 (.IN_OBUF(m0_coef_wdata_dup_0[22]),.OUT_OBUF(m0_coef_wdata[22]));

	qlOBUF QL_INST_F2A_T_12_5 (.IN_OBUF(m0_coef_wdata_dup_0[21]),.OUT_OBUF(m0_coef_wdata[21]));

	qlOBUF QL_INST_F2A_T_12_6 (.IN_OBUF(m0_coef_wdata_dup_0[20]),.OUT_OBUF(m0_coef_wdata[20]));

	qlOBUF QL_INST_F2A_T_12_7 (.IN_OBUF(m0_coef_wdata_dup_0[19]),.OUT_OBUF(m0_coef_wdata[19]));

	qlOBUF QL_INST_F2A_T_12_8 (.IN_OBUF(m0_coef_wdata_dup_0[18]),.OUT_OBUF(m0_coef_wdata[18]));

	qlOBUF QL_INST_F2A_T_12_9 (.IN_OBUF(m0_coef_wdata_dup_0[17]),.OUT_OBUF(m0_coef_wdata[17]));

	qlOBUF QL_INST_F2A_T_12_10 (.IN_OBUF(m0_coef_wdata_dup_0[16]),.OUT_OBUF(m0_coef_wdata[16]));

	qlOBUF QL_INST_F2A_T_12_11 (.IN_OBUF(m0_coef_wdata_dup_0[15]),.OUT_OBUF(m0_coef_wdata[15]));

	qlOBUF QL_INST_F2A_T_12_12 (.IN_OBUF(m0_coef_wdata_dup_0[14]),.OUT_OBUF(m0_coef_wdata[14]));

	qlOBUF QL_INST_F2A_T_12_13 (.IN_OBUF(m0_coef_wdata_dup_0[13]),.OUT_OBUF(m0_coef_wdata[13]));

	qlOBUF QL_INST_F2A_T_12_14 (.IN_OBUF(m0_coef_wdata_dup_0[12]),.OUT_OBUF(m0_coef_wdata[12]));

	qlOBUF QL_INST_F2A_T_12_15 (.IN_OBUF(m0_coef_wdata_dup_0[11]),.OUT_OBUF(m0_coef_wdata[11]));

	qlOBUF QL_INST_F2A_T_12_16 (.IN_OBUF(m0_coef_wdata_dup_0[10]),.OUT_OBUF(m0_coef_wdata[10]));

	qlOBUF QL_INST_F2A_T_12_17 (.IN_OBUF(m0_coef_wdata_dup_0[9]),.OUT_OBUF(m0_coef_wdata[9]));

	qlIBUF QL_INST_A2F_T_12_0 (.IN_IBUF(m0_coef_rdata[29]),.OUT_IBUF(m0_coef_rdata_int[29]));

	qlIBUF QL_INST_A2F_T_12_1 (.IN_IBUF(m0_coef_rdata[28]),.OUT_IBUF(m0_coef_rdata_int[28]));

	qlIBUF QL_INST_A2F_T_12_2 (.IN_IBUF(m0_coef_rdata[27]),.OUT_IBUF(m0_coef_rdata_int[27]));

	qlIBUF QL_INST_A2F_T_12_3 (.IN_IBUF(m0_coef_rdata[26]),.OUT_IBUF(m0_coef_rdata_int[26]));

	qlIBUF QL_INST_A2F_T_12_4 (.IN_IBUF(m0_coef_rdata[25]),.OUT_IBUF(m0_coef_rdata_int[25]));

	qlIBUF QL_INST_A2F_T_12_5 (.IN_IBUF(m0_coef_rdata[24]),.OUT_IBUF(m0_coef_rdata_int[24]));

	qlIBUF QL_INST_A2F_T_12_6 (.IN_IBUF(m0_coef_rdata[23]),.OUT_IBUF(m0_coef_rdata_int[23]));

	qlIBUF QL_INST_A2F_T_12_7 (.IN_IBUF(m0_coef_rdata[22]),.OUT_IBUF(m0_coef_rdata_int[22]));

	qlOBUF QL_INST_F2A_T_13_0 (.IN_OBUF(m1_m0_reset_dup_0),.OUT_OBUF(m1_m0_reset));

	qlOBUF QL_INST_F2A_T_13_1 (.IN_OBUF(m0_coef_wdata_dup_0[8]),.OUT_OBUF(m0_coef_wdata[8]));

	qlOBUF QL_INST_F2A_T_13_2 (.IN_OBUF(m0_coef_wdata_dup_0[7]),.OUT_OBUF(m0_coef_wdata[7]));

	qlOBUF QL_INST_F2A_T_13_3 (.IN_OBUF(m0_coef_wdata_dup_0[6]),.OUT_OBUF(m0_coef_wdata[6]));

	qlOBUF QL_INST_F2A_T_13_4 (.IN_OBUF(m0_coef_wdata_dup_0[5]),.OUT_OBUF(m0_coef_wdata[5]));

	qlOBUF QL_INST_F2A_T_13_5 (.IN_OBUF(m0_coef_wdata_dup_0[4]),.OUT_OBUF(m0_coef_wdata[4]));

	qlOBUF QL_INST_F2A_T_13_6 (.IN_OBUF(m0_coef_wdata_dup_0[3]),.OUT_OBUF(m0_coef_wdata[3]));

	qlOBUF QL_INST_F2A_T_13_7 (.IN_OBUF(m0_coef_wdata_dup_0[2]),.OUT_OBUF(m0_coef_wdata[2]));

	qlOBUF QL_INST_F2A_T_13_8 (.IN_OBUF(m0_coef_wdata_dup_0[1]),.OUT_OBUF(m0_coef_wdata[1]));

	qlOBUF QL_INST_F2A_T_13_9 (.IN_OBUF(m0_coef_wdata_dup_0[0]),.OUT_OBUF(m0_coef_wdata[0]));

	qlOBUF QL_INST_F2A_T_13_10 (.IN_OBUF(m0_coef_waddr_dup_0[11]),.OUT_OBUF(m0_coef_waddr[11]));

	qlOBUF QL_INST_F2A_T_13_11 (.IN_OBUF(m0_coef_waddr_dup_0[10]),.OUT_OBUF(m0_coef_waddr[10]));

	DBUF QL_INST_F2Adef_T_13_0 (.IN_DBUF(GND),.OUT_DBUF(m1_oper0_powerdn));

	qlIBUF QL_INST_A2F_T_13_0 (.IN_IBUF(m0_coef_rdata[21]),.OUT_IBUF(m0_coef_rdata_int[21]));

	qlIBUF QL_INST_A2F_T_13_1 (.IN_IBUF(m0_coef_rdata[20]),.OUT_IBUF(m0_coef_rdata_int[20]));

	qlIBUF QL_INST_A2F_T_13_2 (.IN_IBUF(m0_coef_rdata[19]),.OUT_IBUF(m0_coef_rdata_int[19]));

	qlIBUF QL_INST_A2F_T_13_3 (.IN_IBUF(m0_coef_rdata[18]),.OUT_IBUF(m0_coef_rdata_int[18]));

	qlIBUF QL_INST_A2F_T_13_4 (.IN_IBUF(m0_coef_rdata[17]),.OUT_IBUF(m0_coef_rdata_int[17]));

	qlIBUF QL_INST_A2F_T_13_5 (.IN_IBUF(m0_coef_rdata[16]),.OUT_IBUF(m0_coef_rdata_int[16]));

	qlOBUF QL_INST_F2A_T_14_0 (.IN_OBUF(m0_coef_waddr_dup_0[9]),.OUT_OBUF(m0_coef_waddr[9]));

	qlOBUF QL_INST_F2A_T_14_1 (.IN_OBUF(m0_coef_waddr_dup_0[8]),.OUT_OBUF(m0_coef_waddr[8]));

	qlOBUF QL_INST_F2A_T_14_2 (.IN_OBUF(m0_coef_waddr_dup_0[7]),.OUT_OBUF(m0_coef_waddr[7]));

	qlOBUF QL_INST_F2A_T_14_3 (.IN_OBUF(m0_coef_waddr_dup_0[6]),.OUT_OBUF(m0_coef_waddr[6]));

	qlOBUF QL_INST_F2A_T_14_4 (.IN_OBUF(m0_coef_waddr_dup_0[5]),.OUT_OBUF(m0_coef_waddr[5]));

	qlOBUF QL_INST_F2A_T_14_5 (.IN_OBUF(m0_coef_waddr_dup_0[4]),.OUT_OBUF(m0_coef_waddr[4]));

	qlOBUF QL_INST_F2A_T_14_6 (.IN_OBUF(m0_coef_waddr_dup_0[3]),.OUT_OBUF(m0_coef_waddr[3]));

	qlOBUF QL_INST_F2A_T_14_7 (.IN_OBUF(m0_coef_waddr_dup_0[2]),.OUT_OBUF(m0_coef_waddr[2]));

	qlOBUF QL_INST_F2A_T_14_8 (.IN_OBUF(m0_coef_waddr_dup_0[1]),.OUT_OBUF(m0_coef_waddr[1]));

	qlOBUF QL_INST_F2A_T_14_9 (.IN_OBUF(m0_coef_waddr_dup_0[0]),.OUT_OBUF(m0_coef_waddr[0]));

	qlOBUF QL_INST_F2A_T_14_10 (.IN_OBUF(m0_coef_we_dup_0),.OUT_OBUF(m0_coef_we));

	qlOBUF QL_INST_F2A_T_14_11 (.IN_OBUF(m0_m0_clken_dup_0),.OUT_OBUF(m0_m0_clken));

	qlOBUF QL_INST_F2A_T_14_12 (.IN_OBUF(m0_coef_rmode_dup_0[1]),.OUT_OBUF(m0_coef_rmode[1]));

	qlOBUF QL_INST_F2A_T_14_13 (.IN_OBUF(m0_coef_rmode_dup_0[0]),.OUT_OBUF(m0_coef_rmode[0]));

	qlOBUF QL_INST_F2A_T_14_14 (.IN_OBUF(m0_coef_raddr_dup_0[11]),.OUT_OBUF(m0_coef_raddr[11]));

	qlOBUF QL_INST_F2A_T_14_15 (.IN_OBUF(m0_coef_raddr_dup_0[10]),.OUT_OBUF(m0_coef_raddr[10]));

	qlOBUF QL_INST_F2A_T_14_16 (.IN_OBUF(m0_coef_raddr_dup_0[9]),.OUT_OBUF(m0_coef_raddr[9]));

	qlOBUF QL_INST_F2A_T_14_17 (.IN_OBUF(m0_coef_raddr_dup_0[8]),.OUT_OBUF(m0_coef_raddr[8]));

	qlIBUF QL_INST_A2F_T_14_0 (.IN_IBUF(m0_coef_rdata[15]),.OUT_IBUF(m0_coef_rdata_int[15]));

	qlIBUF QL_INST_A2F_T_14_1 (.IN_IBUF(m0_coef_rdata[14]),.OUT_IBUF(m0_coef_rdata_int[14]));

	qlIBUF QL_INST_A2F_T_14_2 (.IN_IBUF(m0_coef_rdata[13]),.OUT_IBUF(m0_coef_rdata_int[13]));

	qlIBUF QL_INST_A2F_T_14_3 (.IN_IBUF(m0_coef_rdata[12]),.OUT_IBUF(m0_coef_rdata_int[12]));

	qlIBUF QL_INST_A2F_T_14_4 (.IN_IBUF(m0_coef_rdata[11]),.OUT_IBUF(m0_coef_rdata_int[11]));

	qlIBUF QL_INST_A2F_T_14_5 (.IN_IBUF(m0_coef_rdata[10]),.OUT_IBUF(m0_coef_rdata_int[10]));

	qlIBUF QL_INST_A2F_T_14_6 (.IN_IBUF(m0_coef_rdata[9]),.OUT_IBUF(m0_coef_rdata_int[9]));

	qlIBUF QL_INST_A2F_T_14_7 (.IN_IBUF(m0_coef_rdata[8]),.OUT_IBUF(m0_coef_rdata_int[8]));

	qlOBUF QL_INST_F2A_T_15_0 (.IN_OBUF(m0_m0_clr_dup_0),.OUT_OBUF(m0_m0_clr));

	qlOBUF QL_INST_F2A_T_15_1 (.IN_OBUF(m0_coef_raddr_dup_0[7]),.OUT_OBUF(m0_coef_raddr[7]));

	qlOBUF QL_INST_F2A_T_15_2 (.IN_OBUF(m0_coef_raddr_dup_0[6]),.OUT_OBUF(m0_coef_raddr[6]));

	qlOBUF QL_INST_F2A_T_15_3 (.IN_OBUF(m0_coef_raddr_dup_0[5]),.OUT_OBUF(m0_coef_raddr[5]));

	qlOBUF QL_INST_F2A_T_15_4 (.IN_OBUF(m0_coef_raddr_dup_0[4]),.OUT_OBUF(m0_coef_raddr[4]));

	qlOBUF QL_INST_F2A_T_15_5 (.IN_OBUF(m0_coef_raddr_dup_0[3]),.OUT_OBUF(m0_coef_raddr[3]));

	qlOBUF QL_INST_F2A_T_15_6 (.IN_OBUF(m0_coef_raddr_dup_0[2]),.OUT_OBUF(m0_coef_raddr[2]));

	qlOBUF QL_INST_F2A_T_15_7 (.IN_OBUF(m0_coef_raddr_dup_0[1]),.OUT_OBUF(m0_coef_raddr[1]));

	qlOBUF QL_INST_F2A_T_15_8 (.IN_OBUF(m0_coef_raddr_dup_0[0]),.OUT_OBUF(m0_coef_raddr[0]));

	qlOBUF QL_INST_F2A_T_15_9 (.IN_OBUF(m0_coef_wmode_dup_0[1]),.OUT_OBUF(m0_coef_wmode[1]));

	qlOBUF QL_INST_F2A_T_15_10 (.IN_OBUF(m0_coef_wmode_dup_0[0]),.OUT_OBUF(m0_coef_wmode[0]));

	qlIBUF QL_INST_A2F_T_15_0 (.IN_IBUF(m0_coef_rdata[7]),.OUT_IBUF(m0_coef_rdata_int[7]));

	qlIBUF QL_INST_A2F_T_15_1 (.IN_IBUF(m0_coef_rdata[6]),.OUT_IBUF(m0_coef_rdata_int[6]));

	qlIBUF QL_INST_A2F_T_15_2 (.IN_IBUF(m0_coef_rdata[5]),.OUT_IBUF(m0_coef_rdata_int[5]));

	qlIBUF QL_INST_A2F_T_15_3 (.IN_IBUF(m0_coef_rdata[4]),.OUT_IBUF(m0_coef_rdata_int[4]));

	qlIBUF QL_INST_A2F_T_15_4 (.IN_IBUF(m0_coef_rdata[3]),.OUT_IBUF(m0_coef_rdata_int[3]));

	qlIBUF QL_INST_A2F_T_15_5 (.IN_IBUF(m0_coef_rdata[2]),.OUT_IBUF(m0_coef_rdata_int[2]));

	qlIBUF QL_INST_A2F_T_16_0 (.IN_IBUF(m0_coef_rdata[1]),.OUT_IBUF(m0_coef_rdata_int[1]));

	qlIBUF QL_INST_A2F_T_16_1 (.IN_IBUF(m0_coef_rdata[0]),.OUT_IBUF(m0_coef_rdata_int[0]));

	qlOBUF QL_INST_F2A_T_18_8 (.IN_OBUF(m0_m1_outsel_dup_0[5]),.OUT_OBUF(m0_m1_outsel[5]));

	qlOBUF QL_INST_F2A_T_18_9 (.IN_OBUF(m0_m1_outsel_dup_0[4]),.OUT_OBUF(m0_m1_outsel[4]));

	qlOBUF QL_INST_F2A_T_18_10 (.IN_OBUF(m0_m1_outsel_dup_0[3]),.OUT_OBUF(m0_m1_outsel[3]));

	qlOBUF QL_INST_F2A_T_18_11 (.IN_OBUF(m0_m1_outsel_dup_0[2]),.OUT_OBUF(m0_m1_outsel[2]));

	qlOBUF QL_INST_F2A_T_18_12 (.IN_OBUF(m0_m1_outsel_dup_0[1]),.OUT_OBUF(m0_m1_outsel[1]));

	qlOBUF QL_INST_F2A_T_18_13 (.IN_OBUF(m0_m1_outsel_dup_0[0]),.OUT_OBUF(m0_m1_outsel[0]));

	qlOBUF QL_INST_F2A_T_18_14 (.IN_OBUF(m1_m0_csel_dup_0),.OUT_OBUF(m1_m0_csel));

	qlOBUF QL_INST_F2A_T_18_15 (.IN_OBUF(m1_m1_clken_dup_0),.OUT_OBUF(m1_m1_clken));

	qlOBUF QL_INST_F2A_T_18_16 (.IN_OBUF(m1_m0_osel_dup_0),.OUT_OBUF(m1_m0_osel));

	qlOBUF QL_INST_F2A_T_18_17 (.IN_OBUF(m0_m1_csel_dup_0),.OUT_OBUF(m0_m1_csel));

	qlIBUF QL_INST_A2F_T_18_0 (.IN_IBUF(m0_m1_dataout[31]),.OUT_IBUF(m0_m1_dataout_int[31]));

	qlIBUF QL_INST_A2F_T_18_1 (.IN_IBUF(m0_m1_dataout[30]),.OUT_IBUF(m0_m1_dataout_int[30]));

	qlIBUF QL_INST_A2F_T_18_2 (.IN_IBUF(m0_m1_dataout[29]),.OUT_IBUF(m0_m1_dataout_int[29]));

	qlIBUF QL_INST_A2F_T_18_3 (.IN_IBUF(m0_m1_dataout[28]),.OUT_IBUF(m0_m1_dataout_int[28]));

	qlIBUF QL_INST_A2F_T_18_4 (.IN_IBUF(m0_m1_dataout[27]),.OUT_IBUF(m0_m1_dataout_int[27]));

	qlIBUF QL_INST_A2F_T_18_5 (.IN_IBUF(m0_m1_dataout[26]),.OUT_IBUF(m0_m1_dataout_int[26]));

	qlIBUF QL_INST_A2F_T_18_6 (.IN_IBUF(m0_m1_dataout[25]),.OUT_IBUF(m0_m1_dataout_int[25]));

	qlIBUF QL_INST_A2F_T_18_7 (.IN_IBUF(m0_m1_dataout[24]),.OUT_IBUF(m0_m1_dataout_int[24]));

	qlOBUF QL_INST_F2A_T_19_0 (.IN_OBUF(tcdm_wen_p0_dup_0),.OUT_OBUF(tcdm_wen_p0));

	qlOBUF QL_INST_F2A_T_19_1 (.IN_OBUF(tcdm_wen_p1_dup_0),.OUT_OBUF(tcdm_wen_p1));

	qlOBUF QL_INST_F2A_T_19_2 (.IN_OBUF(m1_m0_rnd_dup_0),.OUT_OBUF(m1_m0_rnd));

	qlOBUF QL_INST_F2A_T_19_3 (.IN_OBUF(m1_m1_csel_dup_0),.OUT_OBUF(m1_m1_csel));

	qlOBUF QL_INST_F2A_T_19_4 (.IN_OBUF(m0_coef_rdata_int[31]),.OUT_OBUF(m0_m1_coef_in[31]));

	qlOBUF QL_INST_F2A_T_19_5 (.IN_OBUF(m0_coef_rdata_int[30]),.OUT_OBUF(m0_m1_coef_in[30]));

	qlOBUF QL_INST_F2A_T_19_6 (.IN_OBUF(m0_coef_rdata_int[29]),.OUT_OBUF(m0_m1_coef_in[29]));

	qlOBUF QL_INST_F2A_T_19_7 (.IN_OBUF(m0_coef_rdata_int[28]),.OUT_OBUF(m0_m1_coef_in[28]));

	qlOBUF QL_INST_F2A_T_19_8 (.IN_OBUF(m0_coef_rdata_int[27]),.OUT_OBUF(m0_m1_coef_in[27]));

	qlOBUF QL_INST_F2A_T_19_9 (.IN_OBUF(m0_coef_rdata_int[26]),.OUT_OBUF(m0_m1_coef_in[26]));

	qlOBUF QL_INST_F2A_T_19_10 (.IN_OBUF(m0_coef_rdata_int[25]),.OUT_OBUF(m0_m1_coef_in[25]));

	qlOBUF QL_INST_F2A_T_19_11 (.IN_OBUF(m0_coef_rdata_int[24]),.OUT_OBUF(m0_m1_coef_in[24]));

	qlIBUF QL_INST_A2F_T_19_0 (.IN_IBUF(m0_m1_dataout[23]),.OUT_IBUF(m0_m1_dataout_int[23]));

	qlIBUF QL_INST_A2F_T_19_1 (.IN_IBUF(m0_m1_dataout[22]),.OUT_IBUF(m0_m1_dataout_int[22]));

	qlIBUF QL_INST_A2F_T_19_2 (.IN_IBUF(m0_m1_dataout[21]),.OUT_IBUF(m0_m1_dataout_int[21]));

	qlIBUF QL_INST_A2F_T_19_3 (.IN_IBUF(m0_m1_dataout[20]),.OUT_IBUF(m0_m1_dataout_int[20]));

	qlIBUF QL_INST_A2F_T_19_4 (.IN_IBUF(m0_m1_dataout[19]),.OUT_IBUF(m0_m1_dataout_int[19]));

	qlIBUF QL_INST_A2F_T_19_5 (.IN_IBUF(m0_m1_dataout[18]),.OUT_IBUF(m0_m1_dataout_int[18]));

	qlOBUF QL_INST_F2A_T_20_0 (.IN_OBUF(m0_coef_rdata_int[23]),.OUT_OBUF(m0_m1_coef_in[23]));

	qlOBUF QL_INST_F2A_T_20_1 (.IN_OBUF(m0_coef_rdata_int[22]),.OUT_OBUF(m0_m1_coef_in[22]));

	qlOBUF QL_INST_F2A_T_20_2 (.IN_OBUF(m0_coef_rdata_int[21]),.OUT_OBUF(m0_m1_coef_in[21]));

	qlOBUF QL_INST_F2A_T_20_3 (.IN_OBUF(m0_coef_rdata_int[20]),.OUT_OBUF(m0_m1_coef_in[20]));

	qlOBUF QL_INST_F2A_T_20_4 (.IN_OBUF(m0_coef_rdata_int[19]),.OUT_OBUF(m0_m1_coef_in[19]));

	qlOBUF QL_INST_F2A_T_20_5 (.IN_OBUF(m0_coef_rdata_int[18]),.OUT_OBUF(m0_m1_coef_in[18]));

	qlOBUF QL_INST_F2A_T_20_6 (.IN_OBUF(m0_coef_rdata_int[17]),.OUT_OBUF(m0_m1_coef_in[17]));

	qlOBUF QL_INST_F2A_T_20_7 (.IN_OBUF(m0_coef_rdata_int[16]),.OUT_OBUF(m0_m1_coef_in[16]));

	qlOBUF QL_INST_F2A_T_20_8 (.IN_OBUF(m0_coef_rdata_int[15]),.OUT_OBUF(m0_m1_coef_in[15]));

	qlOBUF QL_INST_F2A_T_20_9 (.IN_OBUF(m0_coef_rdata_int[14]),.OUT_OBUF(m0_m1_coef_in[14]));

	qlOBUF QL_INST_F2A_T_20_10 (.IN_OBUF(m0_coef_rdata_int[13]),.OUT_OBUF(m0_m1_coef_in[13]));

	qlOBUF QL_INST_F2A_T_20_11 (.IN_OBUF(m0_coef_rdata_int[12]),.OUT_OBUF(m0_m1_coef_in[12]));

	qlOBUF QL_INST_F2A_T_20_12 (.IN_OBUF(m0_coef_rdata_int[11]),.OUT_OBUF(m0_m1_coef_in[11]));

	qlOBUF QL_INST_F2A_T_20_13 (.IN_OBUF(m0_coef_rdata_int[10]),.OUT_OBUF(m0_m1_coef_in[10]));

	qlOBUF QL_INST_F2A_T_20_14 (.IN_OBUF(m0_coef_rdata_int[9]),.OUT_OBUF(m0_m1_coef_in[9]));

	qlOBUF QL_INST_F2A_T_20_15 (.IN_OBUF(m0_coef_rdata_int[8]),.OUT_OBUF(m0_m1_coef_in[8]));

	qlOBUF QL_INST_F2A_T_20_16 (.IN_OBUF(m0_coef_rdata_int[7]),.OUT_OBUF(m0_m1_coef_in[7]));

	qlOBUF QL_INST_F2A_T_20_17 (.IN_OBUF(m0_coef_rdata_int[6]),.OUT_OBUF(m0_m1_coef_in[6]));

	qlIBUF QL_INST_A2F_T_20_0 (.IN_IBUF(m0_m1_dataout[17]),.OUT_IBUF(m0_m1_dataout_int[17]));

	qlIBUF QL_INST_A2F_T_20_1 (.IN_IBUF(m0_m1_dataout[16]),.OUT_IBUF(m0_m1_dataout_int[16]));

	qlIBUF QL_INST_A2F_T_20_2 (.IN_IBUF(m0_m1_dataout[15]),.OUT_IBUF(m0_m1_dataout_int[15]));

	qlIBUF QL_INST_A2F_T_20_3 (.IN_IBUF(m0_m1_dataout[14]),.OUT_IBUF(m0_m1_dataout_int[14]));

	qlIBUF QL_INST_A2F_T_20_4 (.IN_IBUF(m0_m1_dataout[13]),.OUT_IBUF(m0_m1_dataout_int[13]));

	qlIBUF QL_INST_A2F_T_20_5 (.IN_IBUF(m0_m1_dataout[12]),.OUT_IBUF(m0_m1_dataout_int[12]));

	qlIBUF QL_INST_A2F_T_20_6 (.IN_IBUF(m0_m1_dataout[11]),.OUT_IBUF(m0_m1_dataout_int[11]));

	qlOBUF QL_INST_F2A_T_21_0 (.IN_OBUF(m0_coef_rdata_int[5]),.OUT_OBUF(m0_m1_coef_in[5]));

	qlOBUF QL_INST_F2A_T_21_1 (.IN_OBUF(m0_coef_rdata_int[4]),.OUT_OBUF(m0_m1_coef_in[4]));

	qlOBUF QL_INST_F2A_T_21_2 (.IN_OBUF(m0_coef_rdata_int[3]),.OUT_OBUF(m0_m1_coef_in[3]));

	qlOBUF QL_INST_F2A_T_21_3 (.IN_OBUF(m0_coef_rdata_int[2]),.OUT_OBUF(m0_m1_coef_in[2]));

	qlOBUF QL_INST_F2A_T_21_4 (.IN_OBUF(m0_coef_rdata_int[1]),.OUT_OBUF(m0_m1_coef_in[1]));

	qlOBUF QL_INST_F2A_T_21_5 (.IN_OBUF(m0_coef_rdata_int[0]),.OUT_OBUF(m0_m1_coef_in[0]));

	qlOBUF QL_INST_F2A_T_21_6 (.IN_OBUF(m0_m1_mode_dup_0[1]),.OUT_OBUF(m0_m1_mode[1]));

	qlOBUF QL_INST_F2A_T_21_7 (.IN_OBUF(m1_m1_osel_dup_0),.OUT_OBUF(m1_m1_osel));

	qlOBUF QL_INST_F2A_T_21_8 (.IN_OBUF(m0_m1_mode_dup_0[0]),.OUT_OBUF(m0_m1_mode[0]));

	qlOBUF QL_INST_F2A_T_21_9 (.IN_OBUF(m0_oper1_rdata_int[31]),.OUT_OBUF(m0_m1_oper_in[31]));

	qlOBUF QL_INST_F2A_T_21_10 (.IN_OBUF(m0_oper1_rdata_int[30]),.OUT_OBUF(m0_m1_oper_in[30]));

	qlOBUF QL_INST_F2A_T_21_11 (.IN_OBUF(m0_oper1_rdata_int[29]),.OUT_OBUF(m0_m1_oper_in[29]));

	qlIBUF QL_INST_A2F_T_21_0 (.IN_IBUF(m0_m1_dataout[10]),.OUT_IBUF(m0_m1_dataout_int[10]));

	qlIBUF QL_INST_A2F_T_21_1 (.IN_IBUF(m0_m1_dataout[9]),.OUT_IBUF(m0_m1_dataout_int[9]));

	qlIBUF QL_INST_A2F_T_21_2 (.IN_IBUF(m0_m1_dataout[8]),.OUT_IBUF(m0_m1_dataout_int[8]));

	qlIBUF QL_INST_A2F_T_21_3 (.IN_IBUF(m0_m1_dataout[7]),.OUT_IBUF(m0_m1_dataout_int[7]));

	qlIBUF QL_INST_A2F_T_21_4 (.IN_IBUF(m0_m1_dataout[6]),.OUT_IBUF(m0_m1_dataout_int[6]));

	qlIBUF QL_INST_A2F_T_21_5 (.IN_IBUF(m0_m1_dataout[5]),.OUT_IBUF(m0_m1_dataout_int[5]));

	qlOBUF QL_INST_F2A_T_22_0 (.IN_OBUF(m0_oper1_rdata_int[28]),.OUT_OBUF(m0_m1_oper_in[28]));

	qlOBUF QL_INST_F2A_T_22_1 (.IN_OBUF(m0_oper1_rdata_int[27]),.OUT_OBUF(m0_m1_oper_in[27]));

	qlOBUF QL_INST_F2A_T_22_2 (.IN_OBUF(m0_oper1_rdata_int[26]),.OUT_OBUF(m0_m1_oper_in[26]));

	qlOBUF QL_INST_F2A_T_22_3 (.IN_OBUF(m0_oper1_rdata_int[25]),.OUT_OBUF(m0_m1_oper_in[25]));

	qlOBUF QL_INST_F2A_T_22_4 (.IN_OBUF(m0_oper1_rdata_int[24]),.OUT_OBUF(m0_m1_oper_in[24]));

	qlOBUF QL_INST_F2A_T_22_5 (.IN_OBUF(m0_oper1_rdata_int[23]),.OUT_OBUF(m0_m1_oper_in[23]));

	qlOBUF QL_INST_F2A_T_22_6 (.IN_OBUF(m0_oper1_rdata_int[22]),.OUT_OBUF(m0_m1_oper_in[22]));

	qlOBUF QL_INST_F2A_T_22_7 (.IN_OBUF(m0_oper1_rdata_int[21]),.OUT_OBUF(m0_m1_oper_in[21]));

	qlOBUF QL_INST_F2A_T_22_8 (.IN_OBUF(m0_oper1_rdata_int[20]),.OUT_OBUF(m0_m1_oper_in[20]));

	qlOBUF QL_INST_F2A_T_22_9 (.IN_OBUF(m0_oper1_rdata_int[19]),.OUT_OBUF(m0_m1_oper_in[19]));

	qlOBUF QL_INST_F2A_T_22_10 (.IN_OBUF(m0_oper1_rdata_int[18]),.OUT_OBUF(m0_m1_oper_in[18]));

	qlOBUF QL_INST_F2A_T_22_11 (.IN_OBUF(m0_oper1_rdata_int[17]),.OUT_OBUF(m0_m1_oper_in[17]));

	qlOBUF QL_INST_F2A_T_22_12 (.IN_OBUF(m0_oper1_rdata_int[16]),.OUT_OBUF(m0_m1_oper_in[16]));

	qlOBUF QL_INST_F2A_T_22_13 (.IN_OBUF(m0_oper1_rdata_int[15]),.OUT_OBUF(m0_m1_oper_in[15]));

	qlOBUF QL_INST_F2A_T_22_14 (.IN_OBUF(m0_oper1_rdata_int[14]),.OUT_OBUF(m0_m1_oper_in[14]));

	qlOBUF QL_INST_F2A_T_22_15 (.IN_OBUF(m0_oper1_rdata_int[13]),.OUT_OBUF(m0_m1_oper_in[13]));

	qlOBUF QL_INST_F2A_T_22_16 (.IN_OBUF(m0_oper1_rdata_int[12]),.OUT_OBUF(m0_m1_oper_in[12]));

	qlOBUF QL_INST_F2A_T_22_17 (.IN_OBUF(m0_oper1_rdata_int[11]),.OUT_OBUF(m0_m1_oper_in[11]));

	qlIBUF QL_INST_A2F_T_22_0 (.IN_IBUF(m0_m1_dataout[4]),.OUT_IBUF(m0_m1_dataout_int[4]));

	qlIBUF QL_INST_A2F_T_22_1 (.IN_IBUF(m0_m1_dataout[3]),.OUT_IBUF(m0_m1_dataout_int[3]));

	qlIBUF QL_INST_A2F_T_22_2 (.IN_IBUF(m0_m1_dataout[2]),.OUT_IBUF(m0_m1_dataout_int[2]));

	qlIBUF QL_INST_A2F_T_22_3 (.IN_IBUF(m0_m1_dataout[1]),.OUT_IBUF(m0_m1_dataout_int[1]));

	qlIBUF QL_INST_A2F_T_22_4 (.IN_IBUF(m0_m1_dataout[0]),.OUT_IBUF(m0_m1_dataout_int[0]));

	qlOBUF QL_INST_F2A_T_23_0 (.IN_OBUF(m0_oper1_rdata_int[10]),.OUT_OBUF(m0_m1_oper_in[10]));

	qlOBUF QL_INST_F2A_T_23_1 (.IN_OBUF(m0_oper1_rdata_int[9]),.OUT_OBUF(m0_m1_oper_in[9]));

	qlOBUF QL_INST_F2A_T_23_2 (.IN_OBUF(m0_oper1_rdata_int[8]),.OUT_OBUF(m0_m1_oper_in[8]));

	qlOBUF QL_INST_F2A_T_23_3 (.IN_OBUF(m0_oper1_rdata_int[7]),.OUT_OBUF(m0_m1_oper_in[7]));

	qlOBUF QL_INST_F2A_T_23_4 (.IN_OBUF(m0_oper1_rdata_int[6]),.OUT_OBUF(m0_m1_oper_in[6]));

	qlOBUF QL_INST_F2A_T_23_5 (.IN_OBUF(m0_oper1_rdata_int[5]),.OUT_OBUF(m0_m1_oper_in[5]));

	qlOBUF QL_INST_F2A_T_23_6 (.IN_OBUF(m0_oper1_rdata_int[4]),.OUT_OBUF(m0_m1_oper_in[4]));

	qlOBUF QL_INST_F2A_T_23_7 (.IN_OBUF(m0_oper1_rdata_int[3]),.OUT_OBUF(m0_m1_oper_in[3]));

	qlOBUF QL_INST_F2A_T_23_8 (.IN_OBUF(m0_oper1_rdata_int[2]),.OUT_OBUF(m0_m1_oper_in[2]));

	qlOBUF QL_INST_F2A_T_23_9 (.IN_OBUF(m0_oper1_rdata_int[1]),.OUT_OBUF(m0_m1_oper_in[1]));

	qlOBUF QL_INST_F2A_T_23_10 (.IN_OBUF(m0_oper1_rdata_int[0]),.OUT_OBUF(m0_m1_oper_in[0]));

	qlOBUF QL_INST_F2A_T_24_16 (.IN_OBUF(m0_oper1_wdata_dup_0[31]),.OUT_OBUF(m0_oper1_wdata[31]));

	qlOBUF QL_INST_F2A_T_24_17 (.IN_OBUF(m0_oper1_wdata_dup_0[30]),.OUT_OBUF(m0_oper1_wdata[30]));

	DBUF QL_INST_F2Adef_T_24_0 (.IN_DBUF(GND),.OUT_DBUF(m0_oper1_powerdn));

	qlOBUF QL_INST_F2A_T_25_0 (.IN_OBUF(m0_oper1_wdata_dup_0[29]),.OUT_OBUF(m0_oper1_wdata[29]));

	qlOBUF QL_INST_F2A_T_25_1 (.IN_OBUF(m0_oper1_wdata_dup_0[28]),.OUT_OBUF(m0_oper1_wdata[28]));

	qlOBUF QL_INST_F2A_T_25_2 (.IN_OBUF(m0_oper1_wdata_dup_0[27]),.OUT_OBUF(m0_oper1_wdata[27]));

	qlOBUF QL_INST_F2A_T_25_3 (.IN_OBUF(m0_oper1_wdata_dup_0[26]),.OUT_OBUF(m0_oper1_wdata[26]));

	qlOBUF QL_INST_F2A_T_25_4 (.IN_OBUF(m0_oper1_wdata_dup_0[25]),.OUT_OBUF(m0_oper1_wdata[25]));

	qlOBUF QL_INST_F2A_T_25_5 (.IN_OBUF(m0_oper1_wdata_dup_0[24]),.OUT_OBUF(m0_oper1_wdata[24]));

	qlOBUF QL_INST_F2A_T_25_6 (.IN_OBUF(m0_oper1_wdata_dup_0[23]),.OUT_OBUF(m0_oper1_wdata[23]));

	qlOBUF QL_INST_F2A_T_25_7 (.IN_OBUF(m0_oper1_wdata_dup_0[22]),.OUT_OBUF(m0_oper1_wdata[22]));

	qlOBUF QL_INST_F2A_T_25_8 (.IN_OBUF(m0_oper1_wdata_dup_0[21]),.OUT_OBUF(m0_oper1_wdata[21]));

	qlOBUF QL_INST_F2A_T_25_9 (.IN_OBUF(m0_oper1_wdata_dup_0[20]),.OUT_OBUF(m0_oper1_wdata[20]));

	qlOBUF QL_INST_F2A_T_25_10 (.IN_OBUF(m0_oper1_wdata_dup_0[19]),.OUT_OBUF(m0_oper1_wdata[19]));

	qlOBUF QL_INST_F2A_T_25_11 (.IN_OBUF(m0_oper1_wdata_dup_0[18]),.OUT_OBUF(m0_oper1_wdata[18]));

	qlIBUF QL_INST_A2F_T_25_1 (.IN_IBUF(m0_oper1_rdata[31]),.OUT_IBUF(m0_oper1_rdata_int[31]));

	qlIBUF QL_INST_A2F_T_25_2 (.IN_IBUF(m0_oper1_rdata[30]),.OUT_IBUF(m0_oper1_rdata_int[30]));

	qlIBUF QL_INST_A2F_T_25_3 (.IN_IBUF(m0_oper1_rdata[29]),.OUT_IBUF(m0_oper1_rdata_int[29]));

	qlIBUF QL_INST_A2F_T_25_4 (.IN_IBUF(m0_oper1_rdata[28]),.OUT_IBUF(m0_oper1_rdata_int[28]));

	qlIBUF QL_INST_A2F_T_25_5 (.IN_IBUF(m0_oper1_rdata[27]),.OUT_IBUF(m0_oper1_rdata_int[27]));

	qlOBUF QL_INST_F2A_T_26_0 (.IN_OBUF(m0_oper1_wdata_dup_0[17]),.OUT_OBUF(m0_oper1_wdata[17]));

	qlOBUF QL_INST_F2A_T_26_1 (.IN_OBUF(m0_oper1_wdata_dup_0[16]),.OUT_OBUF(m0_oper1_wdata[16]));

	qlOBUF QL_INST_F2A_T_26_2 (.IN_OBUF(m0_oper1_wdata_dup_0[15]),.OUT_OBUF(m0_oper1_wdata[15]));

	qlOBUF QL_INST_F2A_T_26_3 (.IN_OBUF(m0_oper1_wdata_dup_0[14]),.OUT_OBUF(m0_oper1_wdata[14]));

	qlOBUF QL_INST_F2A_T_26_4 (.IN_OBUF(m0_oper1_wdata_dup_0[13]),.OUT_OBUF(m0_oper1_wdata[13]));

	qlOBUF QL_INST_F2A_T_26_5 (.IN_OBUF(m0_oper1_wdata_dup_0[12]),.OUT_OBUF(m0_oper1_wdata[12]));

	qlOBUF QL_INST_F2A_T_26_6 (.IN_OBUF(m0_oper1_wdata_dup_0[11]),.OUT_OBUF(m0_oper1_wdata[11]));

	qlOBUF QL_INST_F2A_T_26_7 (.IN_OBUF(m0_oper1_wdata_dup_0[10]),.OUT_OBUF(m0_oper1_wdata[10]));

	qlOBUF QL_INST_F2A_T_26_8 (.IN_OBUF(m0_oper1_wdata_dup_0[9]),.OUT_OBUF(m0_oper1_wdata[9]));

	qlOBUF QL_INST_F2A_T_26_9 (.IN_OBUF(m0_oper1_wdata_dup_0[8]),.OUT_OBUF(m0_oper1_wdata[8]));

	qlOBUF QL_INST_F2A_T_26_10 (.IN_OBUF(m0_oper1_wdata_dup_0[7]),.OUT_OBUF(m0_oper1_wdata[7]));

	qlOBUF QL_INST_F2A_T_26_11 (.IN_OBUF(m0_oper1_wdata_dup_0[6]),.OUT_OBUF(m0_oper1_wdata[6]));

	qlOBUF QL_INST_F2A_T_26_12 (.IN_OBUF(m0_oper1_wdata_dup_0[5]),.OUT_OBUF(m0_oper1_wdata[5]));

	qlOBUF QL_INST_F2A_T_26_13 (.IN_OBUF(m0_oper1_wdata_dup_0[4]),.OUT_OBUF(m0_oper1_wdata[4]));

	qlOBUF QL_INST_F2A_T_26_14 (.IN_OBUF(m0_oper1_wdata_dup_0[3]),.OUT_OBUF(m0_oper1_wdata[3]));

	qlOBUF QL_INST_F2A_T_26_15 (.IN_OBUF(m0_oper1_wdata_dup_0[2]),.OUT_OBUF(m0_oper1_wdata[2]));

	qlOBUF QL_INST_F2A_T_26_16 (.IN_OBUF(m0_oper1_wdata_dup_0[1]),.OUT_OBUF(m0_oper1_wdata[1]));

	qlOBUF QL_INST_F2A_T_26_17 (.IN_OBUF(m0_oper1_wdata_dup_0[0]),.OUT_OBUF(m0_oper1_wdata[0]));

	qlIBUF QL_INST_A2F_T_26_0 (.IN_IBUF(m0_oper1_rdata[26]),.OUT_IBUF(m0_oper1_rdata_int[26]));

	qlIBUF QL_INST_A2F_T_26_1 (.IN_IBUF(m0_oper1_rdata[25]),.OUT_IBUF(m0_oper1_rdata_int[25]));

	qlIBUF QL_INST_A2F_T_26_2 (.IN_IBUF(m0_oper1_rdata[24]),.OUT_IBUF(m0_oper1_rdata_int[24]));

	qlIBUF QL_INST_A2F_T_26_3 (.IN_IBUF(m0_oper1_rdata[23]),.OUT_IBUF(m0_oper1_rdata_int[23]));

	qlIBUF QL_INST_A2F_T_26_4 (.IN_IBUF(m0_oper1_rdata[22]),.OUT_IBUF(m0_oper1_rdata_int[22]));

	qlIBUF QL_INST_A2F_T_26_5 (.IN_IBUF(m0_oper1_rdata[21]),.OUT_IBUF(m0_oper1_rdata_int[21]));

	qlIBUF QL_INST_A2F_T_26_6 (.IN_IBUF(m0_oper1_rdata[20]),.OUT_IBUF(m0_oper1_rdata_int[20]));

	qlIBUF QL_INST_A2F_T_26_7 (.IN_IBUF(m0_oper1_rdata[19]),.OUT_IBUF(m0_oper1_rdata_int[19]));

	qlOBUF QL_INST_F2A_T_27_0 (.IN_OBUF(m0_oper1_waddr_dup_0[11]),.OUT_OBUF(m0_oper1_waddr[11]));

	qlOBUF QL_INST_F2A_T_27_1 (.IN_OBUF(m0_oper1_waddr_dup_0[10]),.OUT_OBUF(m0_oper1_waddr[10]));

	qlOBUF QL_INST_F2A_T_27_2 (.IN_OBUF(m0_oper1_waddr_dup_0[9]),.OUT_OBUF(m0_oper1_waddr[9]));

	qlOBUF QL_INST_F2A_T_27_3 (.IN_OBUF(m0_oper1_waddr_dup_0[8]),.OUT_OBUF(m0_oper1_waddr[8]));

	qlOBUF QL_INST_F2A_T_27_4 (.IN_OBUF(m0_oper1_waddr_dup_0[7]),.OUT_OBUF(m0_oper1_waddr[7]));

	qlOBUF QL_INST_F2A_T_27_5 (.IN_OBUF(m0_oper1_waddr_dup_0[6]),.OUT_OBUF(m0_oper1_waddr[6]));

	qlOBUF QL_INST_F2A_T_27_6 (.IN_OBUF(m0_oper1_waddr_dup_0[5]),.OUT_OBUF(m0_oper1_waddr[5]));

	qlOBUF QL_INST_F2A_T_27_7 (.IN_OBUF(m0_oper1_waddr_dup_0[4]),.OUT_OBUF(m0_oper1_waddr[4]));

	qlOBUF QL_INST_F2A_T_27_8 (.IN_OBUF(m0_oper1_waddr_dup_0[3]),.OUT_OBUF(m0_oper1_waddr[3]));

	qlOBUF QL_INST_F2A_T_27_9 (.IN_OBUF(m0_oper1_waddr_dup_0[2]),.OUT_OBUF(m0_oper1_waddr[2]));

	qlOBUF QL_INST_F2A_T_27_10 (.IN_OBUF(m0_oper1_waddr_dup_0[1]),.OUT_OBUF(m0_oper1_waddr[1]));

	qlOBUF QL_INST_F2A_T_27_11 (.IN_OBUF(m0_oper1_waddr_dup_0[0]),.OUT_OBUF(m0_oper1_waddr[0]));

	qlIBUF QL_INST_A2F_T_27_0 (.IN_IBUF(m0_oper1_rdata[18]),.OUT_IBUF(m0_oper1_rdata_int[18]));

	qlIBUF QL_INST_A2F_T_27_1 (.IN_IBUF(m0_oper1_rdata[17]),.OUT_IBUF(m0_oper1_rdata_int[17]));

	qlIBUF QL_INST_A2F_T_27_2 (.IN_IBUF(m0_oper1_rdata[16]),.OUT_IBUF(m0_oper1_rdata_int[16]));

	qlIBUF QL_INST_A2F_T_27_3 (.IN_IBUF(m0_oper1_rdata[15]),.OUT_IBUF(m0_oper1_rdata_int[15]));

	qlIBUF QL_INST_A2F_T_27_4 (.IN_IBUF(m0_oper1_rdata[14]),.OUT_IBUF(m0_oper1_rdata_int[14]));

	qlIBUF QL_INST_A2F_T_27_5 (.IN_IBUF(m0_oper1_rdata[13]),.OUT_IBUF(m0_oper1_rdata_int[13]));

	qlOBUF QL_INST_F2A_T_28_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_28_padClk),.OUT_OBUF(m1_coef_rclk));

	qlOBUF QL_INST_F2A_T_28_1 (.IN_OBUF(m0_oper1_wmode_dup_0[1]),.OUT_OBUF(m0_oper1_wmode[1]));

	qlOBUF QL_INST_F2A_T_28_2 (.IN_OBUF(m0_oper1_wmode_dup_0[0]),.OUT_OBUF(m0_oper1_wmode[0]));

	qlOBUF QL_INST_F2A_T_28_3 (.IN_OBUF(m0_oper1_raddr_dup_0[11]),.OUT_OBUF(m0_oper1_raddr[11]));

	qlOBUF QL_INST_F2A_T_28_4 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_28_padClk),.OUT_OBUF(m0_m1_clk));

	qlOBUF QL_INST_F2A_T_28_15 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_28_padClk),.OUT_OBUF(m1_oper1_wclk));

	qlOBUF QL_INST_F2A_T_28_16 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_28_padClk),.OUT_OBUF(m0_coef_rclk));

	qlOBUF QL_INST_F2A_T_28_17 (.IN_OBUF(m0_oper1_we_dup_0),.OUT_OBUF(m0_oper1_we));

	qlIBUF QL_INST_A2F_T_28_1 (.IN_IBUF(m0_oper1_rdata[12]),.OUT_IBUF(m0_oper1_rdata_int[12]));

	qlIBUF QL_INST_A2F_T_28_2 (.IN_IBUF(m0_oper1_rdata[11]),.OUT_IBUF(m0_oper1_rdata_int[11]));

	qlIBUF QL_INST_A2F_T_28_3 (.IN_IBUF(m0_oper1_rdata[10]),.OUT_IBUF(m0_oper1_rdata_int[10]));

	qlIBUF QL_INST_A2F_T_28_4 (.IN_IBUF(m0_oper1_rdata[9]),.OUT_IBUF(m0_oper1_rdata_int[9]));

	qlIBUF QL_INST_A2F_T_28_5 (.IN_IBUF(m0_oper1_rdata[8]),.OUT_IBUF(m0_oper1_rdata_int[8]));

	qlIBUF QL_INST_A2F_T_28_6 (.IN_IBUF(m0_oper1_rdata[7]),.OUT_IBUF(m0_oper1_rdata_int[7]));

	qlIBUF QL_INST_A2F_T_28_7 (.IN_IBUF(m0_oper1_rdata[6]),.OUT_IBUF(m0_oper1_rdata_int[6]));

	qlOBUF QL_INST_F2A_T_29_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_29_padClk),.OUT_OBUF(m0_m0_clk));

	qlOBUF QL_INST_F2A_T_29_1 (.IN_OBUF(m0_oper1_raddr_dup_0[10]),.OUT_OBUF(m0_oper1_raddr[10]));

	qlOBUF QL_INST_F2A_T_29_2 (.IN_OBUF(m0_oper1_raddr_dup_0[9]),.OUT_OBUF(m0_oper1_raddr[9]));

	qlOBUF QL_INST_F2A_T_29_3 (.IN_OBUF(m0_oper1_raddr_dup_0[8]),.OUT_OBUF(m0_oper1_raddr[8]));

	qlOBUF QL_INST_F2A_T_29_4 (.IN_OBUF(m0_oper1_raddr_dup_0[7]),.OUT_OBUF(m0_oper1_raddr[7]));

	qlOBUF QL_INST_F2A_T_29_5 (.IN_OBUF(m0_oper1_raddr_dup_0[6]),.OUT_OBUF(m0_oper1_raddr[6]));

	qlOBUF QL_INST_F2A_T_29_6 (.IN_OBUF(m0_oper1_raddr_dup_0[5]),.OUT_OBUF(m0_oper1_raddr[5]));

	qlOBUF QL_INST_F2A_T_29_7 (.IN_OBUF(m0_oper1_raddr_dup_0[4]),.OUT_OBUF(m0_oper1_raddr[4]));

	qlOBUF QL_INST_F2A_T_29_8 (.IN_OBUF(m0_oper1_raddr_dup_0[3]),.OUT_OBUF(m0_oper1_raddr[3]));

	qlOBUF QL_INST_F2A_T_29_9 (.IN_OBUF(m0_oper1_raddr_dup_0[2]),.OUT_OBUF(m0_oper1_raddr[2]));

	qlOBUF QL_INST_F2A_T_29_10 (.IN_OBUF(m0_oper1_raddr_dup_0[1]),.OUT_OBUF(m0_oper1_raddr[1]));

	qlOBUF QL_INST_F2A_T_29_11 (.IN_OBUF(m0_oper1_raddr_dup_0[0]),.OUT_OBUF(m0_oper1_raddr[0]));

	qlIBUF QL_INST_A2F_T_29_0 (.IN_IBUF(m0_oper1_rdata[5]),.OUT_IBUF(m0_oper1_rdata_int[5]));

	qlIBUF QL_INST_A2F_T_29_1 (.IN_IBUF(m0_oper1_rdata[4]),.OUT_IBUF(m0_oper1_rdata_int[4]));

	qlIBUF QL_INST_A2F_T_29_2 (.IN_IBUF(m0_oper1_rdata[3]),.OUT_IBUF(m0_oper1_rdata_int[3]));

	qlIBUF QL_INST_A2F_T_29_3 (.IN_IBUF(m0_oper1_rdata[2]),.OUT_IBUF(m0_oper1_rdata_int[2]));

	qlIBUF QL_INST_A2F_T_29_4 (.IN_IBUF(m0_oper1_rdata[1]),.OUT_IBUF(m0_oper1_rdata_int[1]));

	qlIBUF QL_INST_A2F_T_29_5 (.IN_IBUF(m0_oper1_rdata[0]),.OUT_IBUF(m0_oper1_rdata_int[0]));

	qlOBUF QL_INST_F2A_R_3_0 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_33_padClk),.OUT_OBUF(tcdm_clk_p0));

	qlOBUF QL_INST_F2A_R_3_1 (.IN_OBUF(tcdm_req_p0_dup_0),.OUT_OBUF(tcdm_req_p0));

	qlOBUF QL_INST_F2A_R_3_2 (.IN_OBUF(CLK_int_0__CAND0_TRSTR_33_padClk),.OUT_OBUF(m0_oper0_wclk));

	qlOBUF QL_INST_F2A_R_3_3 (.IN_OBUF(tcdm_be_p0_dup_0[0]),.OUT_OBUF(tcdm_be_p0[0]));

	qlOBUF QL_INST_F2A_R_3_4 (.IN_OBUF(tcdm_be_p0_dup_0[1]),.OUT_OBUF(tcdm_be_p0[1]));

	qlOBUF QL_INST_F2A_R_3_5 (.IN_OBUF(tcdm_be_p0_dup_0[2]),.OUT_OBUF(tcdm_be_p0[2]));

	qlOBUF QL_INST_F2A_R_3_6 (.IN_OBUF(tcdm_be_p0_dup_0[3]),.OUT_OBUF(tcdm_be_p0[3]));

	qlOBUF QL_INST_F2A_R_3_8 (.IN_OBUF(tcdm_addr_p0_dup_0[0]),.OUT_OBUF(tcdm_addr_p0[0]));

	qlOBUF QL_INST_F2A_R_3_9 (.IN_OBUF(tcdm_addr_p0_dup_0[1]),.OUT_OBUF(tcdm_addr_p0[1]));

	qlOBUF QL_INST_F2A_R_3_10 (.IN_OBUF(tcdm_addr_p0_dup_0[2]),.OUT_OBUF(tcdm_addr_p0[2]));

	qlOBUF QL_INST_F2A_R_3_11 (.IN_OBUF(tcdm_addr_p0_dup_0[3]),.OUT_OBUF(tcdm_addr_p0[3]));

	qlIBUF QL_INST_A2F_R_3_0 (.IN_IBUF(tcdm_rdata_p0[0]),.OUT_IBUF(tcdm_rdata_p0_int[0]));

	qlIBUF QL_INST_A2F_R_3_1 (.IN_IBUF(tcdm_rdata_p0[1]),.OUT_IBUF(tcdm_rdata_p0_int[1]));

	qlIBUF QL_INST_A2F_R_3_2 (.IN_IBUF(tcdm_rdata_p0[2]),.OUT_IBUF(tcdm_rdata_p0_int[2]));

	qlIBUF QL_INST_A2F_R_3_3 (.IN_IBUF(tcdm_rdata_p0[3]),.OUT_IBUF(tcdm_rdata_p0_int[3]));

	qlIBUF QL_INST_A2F_R_3_4 (.IN_IBUF(tcdm_valid_p0),.OUT_IBUF(tcdm_valid_p0_int));

	qlIBUF QL_INST_A2F_R_3_5 (.IN_IBUF(tcdm_gnt_p0),.OUT_IBUF(tcdm_gnt_p0_int));

	qlOBUF QL_INST_F2A_R_4_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[0]),.OUT_OBUF(tcdm_wdata_p0[0]));

	qlOBUF QL_INST_F2A_R_4_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[1]),.OUT_OBUF(tcdm_wdata_p0[1]));

	qlOBUF QL_INST_F2A_R_4_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[2]),.OUT_OBUF(tcdm_wdata_p0[2]));

	qlOBUF QL_INST_F2A_R_4_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[3]),.OUT_OBUF(tcdm_wdata_p0[3]));

	qlOBUF QL_INST_F2A_R_4_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[4]),.OUT_OBUF(tcdm_wdata_p0[4]));

	qlOBUF QL_INST_F2A_R_4_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[5]),.OUT_OBUF(tcdm_wdata_p0[5]));

	qlOBUF QL_INST_F2A_R_4_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[6]),.OUT_OBUF(tcdm_wdata_p0[6]));

	qlOBUF QL_INST_F2A_R_4_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[7]),.OUT_OBUF(tcdm_wdata_p0[7]));

	qlOBUF QL_INST_F2A_R_4_9 (.IN_OBUF(tcdm_addr_p0_dup_0[4]),.OUT_OBUF(tcdm_addr_p0[4]));

	qlOBUF QL_INST_F2A_R_4_10 (.IN_OBUF(tcdm_addr_p0_dup_0[5]),.OUT_OBUF(tcdm_addr_p0[5]));

	qlOBUF QL_INST_F2A_R_4_11 (.IN_OBUF(tcdm_addr_p0_dup_0[6]),.OUT_OBUF(tcdm_addr_p0[6]));

	qlOBUF QL_INST_F2A_R_4_12 (.IN_OBUF(tcdm_addr_p0_dup_0[7]),.OUT_OBUF(tcdm_addr_p0[7]));

	qlOBUF QL_INST_F2A_R_4_13 (.IN_OBUF(tcdm_addr_p0_dup_0[8]),.OUT_OBUF(tcdm_addr_p0[8]));

	qlOBUF QL_INST_F2A_R_4_14 (.IN_OBUF(tcdm_addr_p0_dup_0[9]),.OUT_OBUF(tcdm_addr_p0[9]));

	qlIBUF QL_INST_A2F_R_4_0 (.IN_IBUF(tcdm_rdata_p0[4]),.OUT_IBUF(tcdm_rdata_p0_int[4]));

	qlIBUF QL_INST_A2F_R_4_1 (.IN_IBUF(tcdm_rdata_p0[5]),.OUT_IBUF(tcdm_rdata_p0_int[5]));

	qlIBUF QL_INST_A2F_R_4_2 (.IN_IBUF(tcdm_rdata_p0[6]),.OUT_IBUF(tcdm_rdata_p0_int[6]));

	qlIBUF QL_INST_A2F_R_4_3 (.IN_IBUF(tcdm_rdata_p0[7]),.OUT_IBUF(tcdm_rdata_p0_int[7]));

	qlIBUF QL_INST_A2F_R_4_4 (.IN_IBUF(tcdm_rdata_p0[8]),.OUT_IBUF(tcdm_rdata_p0_int[8]));

	qlIBUF QL_INST_A2F_R_4_5 (.IN_IBUF(tcdm_rdata_p0[9]),.OUT_IBUF(tcdm_rdata_p0_int[9]));

	qlIBUF QL_INST_A2F_R_4_6 (.IN_IBUF(tcdm_rdata_p0[10]),.OUT_IBUF(tcdm_rdata_p0_int[10]));

	qlIBUF QL_INST_A2F_R_4_7 (.IN_IBUF(tcdm_rdata_p0[11]),.OUT_IBUF(tcdm_rdata_p0_int[11]));

	qlOBUF QL_INST_F2A_R_5_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[8]),.OUT_OBUF(tcdm_wdata_p0[8]));

	qlOBUF QL_INST_F2A_R_5_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[9]),.OUT_OBUF(tcdm_wdata_p0[9]));

	qlOBUF QL_INST_F2A_R_5_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[10]),.OUT_OBUF(tcdm_wdata_p0[10]));

	qlOBUF QL_INST_F2A_R_5_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[11]),.OUT_OBUF(tcdm_wdata_p0[11]));

	qlOBUF QL_INST_F2A_R_5_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[12]),.OUT_OBUF(tcdm_wdata_p0[12]));

	qlOBUF QL_INST_F2A_R_5_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[13]),.OUT_OBUF(tcdm_wdata_p0[13]));

	qlOBUF QL_INST_F2A_R_5_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[14]),.OUT_OBUF(tcdm_wdata_p0[14]));

	qlOBUF QL_INST_F2A_R_5_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[15]),.OUT_OBUF(tcdm_wdata_p0[15]));

	qlOBUF QL_INST_F2A_R_5_8 (.IN_OBUF(tcdm_addr_p0_dup_0[10]),.OUT_OBUF(tcdm_addr_p0[10]));

	qlOBUF QL_INST_F2A_R_5_9 (.IN_OBUF(tcdm_addr_p0_dup_0[11]),.OUT_OBUF(tcdm_addr_p0[11]));

	qlOBUF QL_INST_F2A_R_5_10 (.IN_OBUF(tcdm_addr_p0_dup_0[12]),.OUT_OBUF(tcdm_addr_p0[12]));

	qlOBUF QL_INST_F2A_R_5_11 (.IN_OBUF(tcdm_addr_p0_dup_0[13]),.OUT_OBUF(tcdm_addr_p0[13]));

	qlIBUF QL_INST_A2F_R_5_0 (.IN_IBUF(tcdm_rdata_p0[12]),.OUT_IBUF(tcdm_rdata_p0_int[12]));

	qlIBUF QL_INST_A2F_R_5_1 (.IN_IBUF(tcdm_rdata_p0[13]),.OUT_IBUF(tcdm_rdata_p0_int[13]));

	qlIBUF QL_INST_A2F_R_5_2 (.IN_IBUF(tcdm_rdata_p0[14]),.OUT_IBUF(tcdm_rdata_p0_int[14]));

	qlIBUF QL_INST_A2F_R_5_3 (.IN_IBUF(tcdm_rdata_p0[15]),.OUT_IBUF(tcdm_rdata_p0_int[15]));

	qlIBUF QL_INST_A2F_R_5_4 (.IN_IBUF(tcdm_fmo_p0),.OUT_IBUF(tcdm_fmo_p0_int));

	qlOBUF QL_INST_F2A_R_6_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[16]),.OUT_OBUF(tcdm_wdata_p0[16]));

	qlOBUF QL_INST_F2A_R_6_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[17]),.OUT_OBUF(tcdm_wdata_p0[17]));

	qlOBUF QL_INST_F2A_R_6_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[18]),.OUT_OBUF(tcdm_wdata_p0[18]));

	qlOBUF QL_INST_F2A_R_6_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[19]),.OUT_OBUF(tcdm_wdata_p0[19]));

	qlOBUF QL_INST_F2A_R_6_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[20]),.OUT_OBUF(tcdm_wdata_p0[20]));

	qlOBUF QL_INST_F2A_R_6_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[21]),.OUT_OBUF(tcdm_wdata_p0[21]));

	qlOBUF QL_INST_F2A_R_6_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[22]),.OUT_OBUF(tcdm_wdata_p0[22]));

	qlOBUF QL_INST_F2A_R_6_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[23]),.OUT_OBUF(tcdm_wdata_p0[23]));

	qlOBUF QL_INST_F2A_R_6_12 (.IN_OBUF(tcdm_addr_p0_dup_0[14]),.OUT_OBUF(tcdm_addr_p0[14]));

	qlOBUF QL_INST_F2A_R_6_13 (.IN_OBUF(tcdm_addr_p0_dup_0[15]),.OUT_OBUF(tcdm_addr_p0[15]));

	qlOBUF QL_INST_F2A_R_6_14 (.IN_OBUF(tcdm_addr_p0_dup_0[16]),.OUT_OBUF(tcdm_addr_p0[16]));

	qlOBUF QL_INST_F2A_R_6_15 (.IN_OBUF(tcdm_addr_p0_dup_0[17]),.OUT_OBUF(tcdm_addr_p0[17]));

	qlOBUF QL_INST_F2A_R_6_16 (.IN_OBUF(tcdm_addr_p0_dup_0[18]),.OUT_OBUF(tcdm_addr_p0[18]));

	qlOBUF QL_INST_F2A_R_6_17 (.IN_OBUF(tcdm_addr_p0_dup_0[19]),.OUT_OBUF(tcdm_addr_p0[19]));

	qlIBUF QL_INST_A2F_R_6_0 (.IN_IBUF(RESET[0]),.OUT_IBUF(RESET_int[0]));

	qlIBUF QL_INST_A2F_R_6_1 (.IN_IBUF(tcdm_rdata_p0[16]),.OUT_IBUF(tcdm_rdata_p0_int[16]));

	qlIBUF QL_INST_A2F_R_6_2 (.IN_IBUF(tcdm_rdata_p0[17]),.OUT_IBUF(tcdm_rdata_p0_int[17]));

	qlIBUF QL_INST_A2F_R_6_3 (.IN_IBUF(tcdm_rdata_p0[18]),.OUT_IBUF(tcdm_rdata_p0_int[18]));

	qlIBUF QL_INST_A2F_R_6_4 (.IN_IBUF(tcdm_rdata_p0[19]),.OUT_IBUF(tcdm_rdata_p0_int[19]));

	qlIBUF QL_INST_A2F_R_6_5 (.IN_IBUF(tcdm_rdata_p0[20]),.OUT_IBUF(tcdm_rdata_p0_int[20]));

	qlIBUF QL_INST_A2F_R_6_6 (.IN_IBUF(tcdm_rdata_p0[21]),.OUT_IBUF(tcdm_rdata_p0_int[21]));

	qlOBUF QL_INST_F2A_R_7_0 (.IN_OBUF(tcdm_wdata_p0_dup_0[24]),.OUT_OBUF(tcdm_wdata_p0[24]));

	qlOBUF QL_INST_F2A_R_7_1 (.IN_OBUF(tcdm_wdata_p0_dup_0[25]),.OUT_OBUF(tcdm_wdata_p0[25]));

	qlOBUF QL_INST_F2A_R_7_2 (.IN_OBUF(tcdm_wdata_p0_dup_0[26]),.OUT_OBUF(tcdm_wdata_p0[26]));

	qlOBUF QL_INST_F2A_R_7_3 (.IN_OBUF(tcdm_wdata_p0_dup_0[27]),.OUT_OBUF(tcdm_wdata_p0[27]));

	qlOBUF QL_INST_F2A_R_7_4 (.IN_OBUF(tcdm_wdata_p0_dup_0[28]),.OUT_OBUF(tcdm_wdata_p0[28]));

	qlOBUF QL_INST_F2A_R_7_5 (.IN_OBUF(tcdm_wdata_p0_dup_0[29]),.OUT_OBUF(tcdm_wdata_p0[29]));

	qlOBUF QL_INST_F2A_R_7_6 (.IN_OBUF(tcdm_wdata_p0_dup_0[30]),.OUT_OBUF(tcdm_wdata_p0[30]));

	qlOBUF QL_INST_F2A_R_7_7 (.IN_OBUF(tcdm_wdata_p0_dup_0[31]),.OUT_OBUF(tcdm_wdata_p0[31]));

	qlIBUF QL_INST_A2F_R_7_0 (.IN_IBUF(tcdm_rdata_p0[22]),.OUT_IBUF(tcdm_rdata_p0_int[22]));

	qlIBUF QL_INST_A2F_R_7_1 (.IN_IBUF(tcdm_rdata_p0[23]),.OUT_IBUF(tcdm_rdata_p0_int[23]));

	qlIBUF QL_INST_A2F_R_7_2 (.IN_IBUF(tcdm_rdata_p0[24]),.OUT_IBUF(tcdm_rdata_p0_int[24]));

	qlIBUF QL_INST_A2F_R_7_3 (.IN_IBUF(tcdm_rdata_p0[25]),.OUT_IBUF(tcdm_rdata_p0_int[25]));

	qlIBUF QL_INST_A2F_R_7_4 (.IN_IBUF(tcdm_rdata_p0[26]),.OUT_IBUF(tcdm_rdata_p0_int[26]));

	qlIBUF QL_INST_A2F_R_7_5 (.IN_IBUF(tcdm_rdata_p0[27]),.OUT_IBUF(tcdm_rdata_p0_int[27]));

	qlIBUF QL_INST_A2F_R_8_0 (.IN_IBUF(tcdm_rdata_p0[28]),.OUT_IBUF(tcdm_rdata_p0_int[28]));

	qlIBUF QL_INST_A2F_R_8_1 (.IN_IBUF(tcdm_rdata_p0[29]),.OUT_IBUF(tcdm_rdata_p0_int[29]));

	qlIBUF QL_INST_A2F_R_8_2 (.IN_IBUF(tcdm_rdata_p0[30]),.OUT_IBUF(tcdm_rdata_p0_int[30]));

	qlIBUF QL_INST_A2F_R_8_3 (.IN_IBUF(tcdm_rdata_p0[31]),.OUT_IBUF(tcdm_rdata_p0_int[31]));

	qlOBUF QL_INST_F2A_R_9_0 (.IN_OBUF(CLK_int_0__CAND0_TRSBR_33_padClk),.OUT_OBUF(tcdm_clk_p1));

	qlOBUF QL_INST_F2A_R_9_1 (.IN_OBUF(tcdm_req_p1_dup_0),.OUT_OBUF(tcdm_req_p1));

	qlOBUF QL_INST_F2A_R_9_2 (.IN_OBUF(m0_m0_sat_dup_0),.OUT_OBUF(m0_m0_sat));

	qlOBUF QL_INST_F2A_R_9_3 (.IN_OBUF(tcdm_be_p1_dup_0[0]),.OUT_OBUF(tcdm_be_p1[0]));

	qlOBUF QL_INST_F2A_R_9_4 (.IN_OBUF(tcdm_be_p1_dup_0[1]),.OUT_OBUF(tcdm_be_p1[1]));

	qlOBUF QL_INST_F2A_R_9_5 (.IN_OBUF(tcdm_be_p1_dup_0[2]),.OUT_OBUF(tcdm_be_p1[2]));

	qlOBUF QL_INST_F2A_R_9_6 (.IN_OBUF(tcdm_be_p1_dup_0[3]),.OUT_OBUF(tcdm_be_p1[3]));

	qlOBUF QL_INST_F2A_R_9_8 (.IN_OBUF(tcdm_addr_p1_dup_0[0]),.OUT_OBUF(tcdm_addr_p1[0]));

	qlOBUF QL_INST_F2A_R_9_9 (.IN_OBUF(tcdm_addr_p1_dup_0[1]),.OUT_OBUF(tcdm_addr_p1[1]));

	qlOBUF QL_INST_F2A_R_9_10 (.IN_OBUF(tcdm_addr_p1_dup_0[2]),.OUT_OBUF(tcdm_addr_p1[2]));

	qlOBUF QL_INST_F2A_R_9_11 (.IN_OBUF(tcdm_addr_p1_dup_0[3]),.OUT_OBUF(tcdm_addr_p1[3]));

	qlIBUF QL_INST_A2F_R_9_0 (.IN_IBUF(tcdm_rdata_p1[0]),.OUT_IBUF(tcdm_rdata_p1_int[0]));

	qlIBUF QL_INST_A2F_R_9_1 (.IN_IBUF(tcdm_rdata_p1[1]),.OUT_IBUF(tcdm_rdata_p1_int[1]));

	qlIBUF QL_INST_A2F_R_9_2 (.IN_IBUF(tcdm_rdata_p1[2]),.OUT_IBUF(tcdm_rdata_p1_int[2]));

	qlIBUF QL_INST_A2F_R_9_3 (.IN_IBUF(tcdm_rdata_p1[3]),.OUT_IBUF(tcdm_rdata_p1_int[3]));

	qlIBUF QL_INST_A2F_R_9_4 (.IN_IBUF(tcdm_valid_p1),.OUT_IBUF(tcdm_valid_p1_int));

	qlIBUF QL_INST_A2F_R_9_5 (.IN_IBUF(tcdm_gnt_p1),.OUT_IBUF(tcdm_gnt_p1_int));

	qlOBUF QL_INST_F2A_R_10_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[0]),.OUT_OBUF(tcdm_wdata_p1[0]));

	qlOBUF QL_INST_F2A_R_10_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[1]),.OUT_OBUF(tcdm_wdata_p1[1]));

	qlOBUF QL_INST_F2A_R_10_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[2]),.OUT_OBUF(tcdm_wdata_p1[2]));

	qlOBUF QL_INST_F2A_R_10_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[3]),.OUT_OBUF(tcdm_wdata_p1[3]));

	qlOBUF QL_INST_F2A_R_10_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[4]),.OUT_OBUF(tcdm_wdata_p1[4]));

	qlOBUF QL_INST_F2A_R_10_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[5]),.OUT_OBUF(tcdm_wdata_p1[5]));

	qlOBUF QL_INST_F2A_R_10_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[6]),.OUT_OBUF(tcdm_wdata_p1[6]));

	qlOBUF QL_INST_F2A_R_10_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[7]),.OUT_OBUF(tcdm_wdata_p1[7]));

	qlOBUF QL_INST_F2A_R_10_9 (.IN_OBUF(tcdm_addr_p1_dup_0[4]),.OUT_OBUF(tcdm_addr_p1[4]));

	qlOBUF QL_INST_F2A_R_10_10 (.IN_OBUF(tcdm_addr_p1_dup_0[5]),.OUT_OBUF(tcdm_addr_p1[5]));

	qlOBUF QL_INST_F2A_R_10_11 (.IN_OBUF(tcdm_addr_p1_dup_0[6]),.OUT_OBUF(tcdm_addr_p1[6]));

	qlOBUF QL_INST_F2A_R_10_12 (.IN_OBUF(tcdm_addr_p1_dup_0[7]),.OUT_OBUF(tcdm_addr_p1[7]));

	qlOBUF QL_INST_F2A_R_10_13 (.IN_OBUF(tcdm_addr_p1_dup_0[8]),.OUT_OBUF(tcdm_addr_p1[8]));

	qlOBUF QL_INST_F2A_R_10_14 (.IN_OBUF(tcdm_addr_p1_dup_0[9]),.OUT_OBUF(tcdm_addr_p1[9]));

	qlIBUF QL_INST_A2F_R_10_0 (.IN_IBUF(tcdm_rdata_p1[4]),.OUT_IBUF(tcdm_rdata_p1_int[4]));

	qlIBUF QL_INST_A2F_R_10_1 (.IN_IBUF(tcdm_rdata_p1[5]),.OUT_IBUF(tcdm_rdata_p1_int[5]));

	qlIBUF QL_INST_A2F_R_10_2 (.IN_IBUF(tcdm_rdata_p1[6]),.OUT_IBUF(tcdm_rdata_p1_int[6]));

	qlIBUF QL_INST_A2F_R_10_3 (.IN_IBUF(tcdm_rdata_p1[7]),.OUT_IBUF(tcdm_rdata_p1_int[7]));

	qlIBUF QL_INST_A2F_R_10_4 (.IN_IBUF(tcdm_rdata_p1[8]),.OUT_IBUF(tcdm_rdata_p1_int[8]));

	qlIBUF QL_INST_A2F_R_10_5 (.IN_IBUF(tcdm_rdata_p1[9]),.OUT_IBUF(tcdm_rdata_p1_int[9]));

	qlIBUF QL_INST_A2F_R_10_6 (.IN_IBUF(tcdm_rdata_p1[10]),.OUT_IBUF(tcdm_rdata_p1_int[10]));

	qlIBUF QL_INST_A2F_R_10_7 (.IN_IBUF(tcdm_rdata_p1[11]),.OUT_IBUF(tcdm_rdata_p1_int[11]));

	qlOBUF QL_INST_F2A_R_11_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[8]),.OUT_OBUF(tcdm_wdata_p1[8]));

	qlOBUF QL_INST_F2A_R_11_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[9]),.OUT_OBUF(tcdm_wdata_p1[9]));

	qlOBUF QL_INST_F2A_R_11_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[10]),.OUT_OBUF(tcdm_wdata_p1[10]));

	qlOBUF QL_INST_F2A_R_11_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[11]),.OUT_OBUF(tcdm_wdata_p1[11]));

	qlOBUF QL_INST_F2A_R_11_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[12]),.OUT_OBUF(tcdm_wdata_p1[12]));

	qlOBUF QL_INST_F2A_R_11_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[13]),.OUT_OBUF(tcdm_wdata_p1[13]));

	qlOBUF QL_INST_F2A_R_11_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[14]),.OUT_OBUF(tcdm_wdata_p1[14]));

	qlOBUF QL_INST_F2A_R_11_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[15]),.OUT_OBUF(tcdm_wdata_p1[15]));

	qlOBUF QL_INST_F2A_R_11_8 (.IN_OBUF(tcdm_addr_p1_dup_0[10]),.OUT_OBUF(tcdm_addr_p1[10]));

	qlOBUF QL_INST_F2A_R_11_9 (.IN_OBUF(tcdm_addr_p1_dup_0[11]),.OUT_OBUF(tcdm_addr_p1[11]));

	qlOBUF QL_INST_F2A_R_11_10 (.IN_OBUF(tcdm_addr_p1_dup_0[12]),.OUT_OBUF(tcdm_addr_p1[12]));

	qlOBUF QL_INST_F2A_R_11_11 (.IN_OBUF(tcdm_addr_p1_dup_0[13]),.OUT_OBUF(tcdm_addr_p1[13]));

	qlIBUF QL_INST_A2F_R_11_0 (.IN_IBUF(tcdm_rdata_p1[12]),.OUT_IBUF(tcdm_rdata_p1_int[12]));

	qlIBUF QL_INST_A2F_R_11_1 (.IN_IBUF(tcdm_rdata_p1[13]),.OUT_IBUF(tcdm_rdata_p1_int[13]));

	qlIBUF QL_INST_A2F_R_11_2 (.IN_IBUF(tcdm_rdata_p1[14]),.OUT_IBUF(tcdm_rdata_p1_int[14]));

	qlIBUF QL_INST_A2F_R_11_3 (.IN_IBUF(tcdm_rdata_p1[15]),.OUT_IBUF(tcdm_rdata_p1_int[15]));

	qlIBUF QL_INST_A2F_R_11_4 (.IN_IBUF(tcdm_fmo_p1),.OUT_IBUF(tcdm_fmo_p1_int));

	qlOBUF QL_INST_F2A_R_12_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[16]),.OUT_OBUF(tcdm_wdata_p1[16]));

	qlOBUF QL_INST_F2A_R_12_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[17]),.OUT_OBUF(tcdm_wdata_p1[17]));

	qlOBUF QL_INST_F2A_R_12_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[18]),.OUT_OBUF(tcdm_wdata_p1[18]));

	qlOBUF QL_INST_F2A_R_12_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[19]),.OUT_OBUF(tcdm_wdata_p1[19]));

	qlOBUF QL_INST_F2A_R_12_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[20]),.OUT_OBUF(tcdm_wdata_p1[20]));

	qlOBUF QL_INST_F2A_R_12_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[21]),.OUT_OBUF(tcdm_wdata_p1[21]));

	qlOBUF QL_INST_F2A_R_12_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[22]),.OUT_OBUF(tcdm_wdata_p1[22]));

	qlOBUF QL_INST_F2A_R_12_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[23]),.OUT_OBUF(tcdm_wdata_p1[23]));

	qlOBUF QL_INST_F2A_R_12_12 (.IN_OBUF(tcdm_addr_p1_dup_0[14]),.OUT_OBUF(tcdm_addr_p1[14]));

	qlOBUF QL_INST_F2A_R_12_13 (.IN_OBUF(tcdm_addr_p1_dup_0[15]),.OUT_OBUF(tcdm_addr_p1[15]));

	qlOBUF QL_INST_F2A_R_12_14 (.IN_OBUF(tcdm_addr_p1_dup_0[16]),.OUT_OBUF(tcdm_addr_p1[16]));

	qlOBUF QL_INST_F2A_R_12_15 (.IN_OBUF(tcdm_addr_p1_dup_0[17]),.OUT_OBUF(tcdm_addr_p1[17]));

	qlOBUF QL_INST_F2A_R_12_16 (.IN_OBUF(tcdm_addr_p1_dup_0[18]),.OUT_OBUF(tcdm_addr_p1[18]));

	qlOBUF QL_INST_F2A_R_12_17 (.IN_OBUF(tcdm_addr_p1_dup_0[19]),.OUT_OBUF(tcdm_addr_p1[19]));

	qlIBUF QL_INST_A2F_R_12_1 (.IN_IBUF(tcdm_rdata_p1[16]),.OUT_IBUF(tcdm_rdata_p1_int[16]));

	qlIBUF QL_INST_A2F_R_12_2 (.IN_IBUF(tcdm_rdata_p1[17]),.OUT_IBUF(tcdm_rdata_p1_int[17]));

	qlIBUF QL_INST_A2F_R_12_3 (.IN_IBUF(tcdm_rdata_p1[18]),.OUT_IBUF(tcdm_rdata_p1_int[18]));

	qlIBUF QL_INST_A2F_R_12_4 (.IN_IBUF(tcdm_rdata_p1[19]),.OUT_IBUF(tcdm_rdata_p1_int[19]));

	qlIBUF QL_INST_A2F_R_12_5 (.IN_IBUF(tcdm_rdata_p1[20]),.OUT_IBUF(tcdm_rdata_p1_int[20]));

	qlIBUF QL_INST_A2F_R_12_6 (.IN_IBUF(tcdm_rdata_p1[21]),.OUT_IBUF(tcdm_rdata_p1_int[21]));

	qlOBUF QL_INST_F2A_R_13_0 (.IN_OBUF(tcdm_wdata_p1_dup_0[24]),.OUT_OBUF(tcdm_wdata_p1[24]));

	qlOBUF QL_INST_F2A_R_13_1 (.IN_OBUF(tcdm_wdata_p1_dup_0[25]),.OUT_OBUF(tcdm_wdata_p1[25]));

	qlOBUF QL_INST_F2A_R_13_2 (.IN_OBUF(tcdm_wdata_p1_dup_0[26]),.OUT_OBUF(tcdm_wdata_p1[26]));

	qlOBUF QL_INST_F2A_R_13_3 (.IN_OBUF(tcdm_wdata_p1_dup_0[27]),.OUT_OBUF(tcdm_wdata_p1[27]));

	qlOBUF QL_INST_F2A_R_13_4 (.IN_OBUF(tcdm_wdata_p1_dup_0[28]),.OUT_OBUF(tcdm_wdata_p1[28]));

	qlOBUF QL_INST_F2A_R_13_5 (.IN_OBUF(tcdm_wdata_p1_dup_0[29]),.OUT_OBUF(tcdm_wdata_p1[29]));

	qlOBUF QL_INST_F2A_R_13_6 (.IN_OBUF(tcdm_wdata_p1_dup_0[30]),.OUT_OBUF(tcdm_wdata_p1[30]));

	qlOBUF QL_INST_F2A_R_13_7 (.IN_OBUF(tcdm_wdata_p1_dup_0[31]),.OUT_OBUF(tcdm_wdata_p1[31]));

	qlIBUF QL_INST_A2F_R_13_0 (.IN_IBUF(tcdm_rdata_p1[22]),.OUT_IBUF(tcdm_rdata_p1_int[22]));

	qlIBUF QL_INST_A2F_R_13_1 (.IN_IBUF(tcdm_rdata_p1[23]),.OUT_IBUF(tcdm_rdata_p1_int[23]));

	qlIBUF QL_INST_A2F_R_13_2 (.IN_IBUF(tcdm_rdata_p1[24]),.OUT_IBUF(tcdm_rdata_p1_int[24]));

	qlIBUF QL_INST_A2F_R_13_3 (.IN_IBUF(tcdm_rdata_p1[25]),.OUT_IBUF(tcdm_rdata_p1_int[25]));

	qlIBUF QL_INST_A2F_R_13_4 (.IN_IBUF(tcdm_rdata_p1[26]),.OUT_IBUF(tcdm_rdata_p1_int[26]));

	qlIBUF QL_INST_A2F_R_13_5 (.IN_IBUF(tcdm_rdata_p1[27]),.OUT_IBUF(tcdm_rdata_p1_int[27]));

	qlIBUF QL_INST_A2F_R_14_0 (.IN_IBUF(tcdm_rdata_p1[28]),.OUT_IBUF(tcdm_rdata_p1_int[28]));

	qlIBUF QL_INST_A2F_R_14_1 (.IN_IBUF(tcdm_rdata_p1[29]),.OUT_IBUF(tcdm_rdata_p1_int[29]));

	qlIBUF QL_INST_A2F_R_14_2 (.IN_IBUF(tcdm_rdata_p1[30]),.OUT_IBUF(tcdm_rdata_p1_int[30]));

	qlIBUF QL_INST_A2F_R_14_3 (.IN_IBUF(tcdm_rdata_p1[31]),.OUT_IBUF(tcdm_rdata_p1_int[31]));

	qlOBUF QL_INST_F2A_R_17_0 (.IN_OBUF(CLK_int_0__CAND0_BRSTR_33_padClk),.OUT_OBUF(tcdm_clk_p2));

	qlOBUF QL_INST_F2A_R_17_1 (.IN_OBUF(tcdm_req_p2_dup_0),.OUT_OBUF(tcdm_req_p2));

	qlOBUF QL_INST_F2A_R_17_2 (.IN_OBUF(m1_m1_rnd_dup_0),.OUT_OBUF(m1_m1_rnd));

	qlOBUF QL_INST_F2A_R_17_3 (.IN_OBUF(tcdm_be_p2_dup_0[0]),.OUT_OBUF(tcdm_be_p2[0]));

	qlOBUF QL_INST_F2A_R_17_4 (.IN_OBUF(tcdm_be_p2_dup_0[1]),.OUT_OBUF(tcdm_be_p2[1]));

	qlOBUF QL_INST_F2A_R_17_5 (.IN_OBUF(tcdm_be_p2_dup_0[2]),.OUT_OBUF(tcdm_be_p2[2]));

	qlOBUF QL_INST_F2A_R_17_6 (.IN_OBUF(tcdm_be_p2_dup_0[3]),.OUT_OBUF(tcdm_be_p2[3]));

	qlOBUF QL_INST_F2A_R_17_8 (.IN_OBUF(tcdm_addr_p2_dup_0[0]),.OUT_OBUF(tcdm_addr_p2[0]));

	qlOBUF QL_INST_F2A_R_17_9 (.IN_OBUF(tcdm_addr_p2_dup_0[1]),.OUT_OBUF(tcdm_addr_p2[1]));

	qlOBUF QL_INST_F2A_R_17_10 (.IN_OBUF(tcdm_addr_p2_dup_0[2]),.OUT_OBUF(tcdm_addr_p2[2]));

	qlOBUF QL_INST_F2A_R_17_11 (.IN_OBUF(tcdm_addr_p2_dup_0[3]),.OUT_OBUF(tcdm_addr_p2[3]));

	qlIBUF QL_INST_A2F_R_17_0 (.IN_IBUF(tcdm_rdata_p2[0]),.OUT_IBUF(tcdm_rdata_p2_int[0]));

	qlIBUF QL_INST_A2F_R_17_1 (.IN_IBUF(tcdm_rdata_p2[1]),.OUT_IBUF(tcdm_rdata_p2_int[1]));

	qlIBUF QL_INST_A2F_R_17_2 (.IN_IBUF(tcdm_rdata_p2[2]),.OUT_IBUF(tcdm_rdata_p2_int[2]));

	qlIBUF QL_INST_A2F_R_17_3 (.IN_IBUF(tcdm_rdata_p2[3]),.OUT_IBUF(tcdm_rdata_p2_int[3]));

	qlIBUF QL_INST_A2F_R_17_4 (.IN_IBUF(tcdm_valid_p2),.OUT_IBUF(tcdm_valid_p2_int));

	qlIBUF QL_INST_A2F_R_17_5 (.IN_IBUF(tcdm_gnt_p2),.OUT_IBUF(tcdm_gnt_p2_int));

	qlOBUF QL_INST_F2A_R_18_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[0]),.OUT_OBUF(tcdm_wdata_p2[0]));

	qlOBUF QL_INST_F2A_R_18_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[1]),.OUT_OBUF(tcdm_wdata_p2[1]));

	qlOBUF QL_INST_F2A_R_18_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[2]),.OUT_OBUF(tcdm_wdata_p2[2]));

	qlOBUF QL_INST_F2A_R_18_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[3]),.OUT_OBUF(tcdm_wdata_p2[3]));

	qlOBUF QL_INST_F2A_R_18_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[4]),.OUT_OBUF(tcdm_wdata_p2[4]));

	qlOBUF QL_INST_F2A_R_18_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[5]),.OUT_OBUF(tcdm_wdata_p2[5]));

	qlOBUF QL_INST_F2A_R_18_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[6]),.OUT_OBUF(tcdm_wdata_p2[6]));

	qlOBUF QL_INST_F2A_R_18_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[7]),.OUT_OBUF(tcdm_wdata_p2[7]));

	qlOBUF QL_INST_F2A_R_18_9 (.IN_OBUF(tcdm_addr_p2_dup_0[4]),.OUT_OBUF(tcdm_addr_p2[4]));

	qlOBUF QL_INST_F2A_R_18_10 (.IN_OBUF(tcdm_addr_p2_dup_0[5]),.OUT_OBUF(tcdm_addr_p2[5]));

	qlOBUF QL_INST_F2A_R_18_11 (.IN_OBUF(tcdm_addr_p2_dup_0[6]),.OUT_OBUF(tcdm_addr_p2[6]));

	qlOBUF QL_INST_F2A_R_18_12 (.IN_OBUF(tcdm_addr_p2_dup_0[7]),.OUT_OBUF(tcdm_addr_p2[7]));

	qlOBUF QL_INST_F2A_R_18_13 (.IN_OBUF(tcdm_addr_p2_dup_0[8]),.OUT_OBUF(tcdm_addr_p2[8]));

	qlOBUF QL_INST_F2A_R_18_14 (.IN_OBUF(tcdm_addr_p2_dup_0[9]),.OUT_OBUF(tcdm_addr_p2[9]));

	qlIBUF QL_INST_A2F_R_18_0 (.IN_IBUF(tcdm_rdata_p2[4]),.OUT_IBUF(tcdm_rdata_p2_int[4]));

	qlIBUF QL_INST_A2F_R_18_1 (.IN_IBUF(tcdm_rdata_p2[5]),.OUT_IBUF(tcdm_rdata_p2_int[5]));

	qlIBUF QL_INST_A2F_R_18_2 (.IN_IBUF(tcdm_rdata_p2[6]),.OUT_IBUF(tcdm_rdata_p2_int[6]));

	qlIBUF QL_INST_A2F_R_18_3 (.IN_IBUF(tcdm_rdata_p2[7]),.OUT_IBUF(tcdm_rdata_p2_int[7]));

	qlIBUF QL_INST_A2F_R_18_4 (.IN_IBUF(tcdm_rdata_p2[8]),.OUT_IBUF(tcdm_rdata_p2_int[8]));

	qlIBUF QL_INST_A2F_R_18_5 (.IN_IBUF(tcdm_rdata_p2[9]),.OUT_IBUF(tcdm_rdata_p2_int[9]));

	qlIBUF QL_INST_A2F_R_18_6 (.IN_IBUF(tcdm_rdata_p2[10]),.OUT_IBUF(tcdm_rdata_p2_int[10]));

	qlIBUF QL_INST_A2F_R_18_7 (.IN_IBUF(tcdm_rdata_p2[11]),.OUT_IBUF(tcdm_rdata_p2_int[11]));

	qlOBUF QL_INST_F2A_R_19_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[8]),.OUT_OBUF(tcdm_wdata_p2[8]));

	qlOBUF QL_INST_F2A_R_19_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[9]),.OUT_OBUF(tcdm_wdata_p2[9]));

	qlOBUF QL_INST_F2A_R_19_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[10]),.OUT_OBUF(tcdm_wdata_p2[10]));

	qlOBUF QL_INST_F2A_R_19_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[11]),.OUT_OBUF(tcdm_wdata_p2[11]));

	qlOBUF QL_INST_F2A_R_19_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[12]),.OUT_OBUF(tcdm_wdata_p2[12]));

	qlOBUF QL_INST_F2A_R_19_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[13]),.OUT_OBUF(tcdm_wdata_p2[13]));

	qlOBUF QL_INST_F2A_R_19_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[14]),.OUT_OBUF(tcdm_wdata_p2[14]));

	qlOBUF QL_INST_F2A_R_19_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[15]),.OUT_OBUF(tcdm_wdata_p2[15]));

	qlOBUF QL_INST_F2A_R_19_8 (.IN_OBUF(tcdm_addr_p2_dup_0[10]),.OUT_OBUF(tcdm_addr_p2[10]));

	qlOBUF QL_INST_F2A_R_19_9 (.IN_OBUF(tcdm_addr_p2_dup_0[11]),.OUT_OBUF(tcdm_addr_p2[11]));

	qlOBUF QL_INST_F2A_R_19_10 (.IN_OBUF(tcdm_addr_p2_dup_0[12]),.OUT_OBUF(tcdm_addr_p2[12]));

	qlOBUF QL_INST_F2A_R_19_11 (.IN_OBUF(tcdm_addr_p2_dup_0[13]),.OUT_OBUF(tcdm_addr_p2[13]));

	qlIBUF QL_INST_A2F_R_19_0 (.IN_IBUF(tcdm_rdata_p2[12]),.OUT_IBUF(tcdm_rdata_p2_int[12]));

	qlIBUF QL_INST_A2F_R_19_1 (.IN_IBUF(tcdm_rdata_p2[13]),.OUT_IBUF(tcdm_rdata_p2_int[13]));

	qlIBUF QL_INST_A2F_R_19_2 (.IN_IBUF(tcdm_rdata_p2[14]),.OUT_IBUF(tcdm_rdata_p2_int[14]));

	qlIBUF QL_INST_A2F_R_19_3 (.IN_IBUF(tcdm_rdata_p2[15]),.OUT_IBUF(tcdm_rdata_p2_int[15]));

	qlIBUF QL_INST_A2F_R_19_4 (.IN_IBUF(tcdm_fmo_p2),.OUT_IBUF(tcdm_fmo_p2_int));

	qlOBUF QL_INST_F2A_R_20_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[16]),.OUT_OBUF(tcdm_wdata_p2[16]));

	qlOBUF QL_INST_F2A_R_20_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[17]),.OUT_OBUF(tcdm_wdata_p2[17]));

	qlOBUF QL_INST_F2A_R_20_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[18]),.OUT_OBUF(tcdm_wdata_p2[18]));

	qlOBUF QL_INST_F2A_R_20_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[19]),.OUT_OBUF(tcdm_wdata_p2[19]));

	qlOBUF QL_INST_F2A_R_20_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[20]),.OUT_OBUF(tcdm_wdata_p2[20]));

	qlOBUF QL_INST_F2A_R_20_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[21]),.OUT_OBUF(tcdm_wdata_p2[21]));

	qlOBUF QL_INST_F2A_R_20_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[22]),.OUT_OBUF(tcdm_wdata_p2[22]));

	qlOBUF QL_INST_F2A_R_20_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[23]),.OUT_OBUF(tcdm_wdata_p2[23]));

	qlOBUF QL_INST_F2A_R_20_12 (.IN_OBUF(tcdm_addr_p2_dup_0[14]),.OUT_OBUF(tcdm_addr_p2[14]));

	qlOBUF QL_INST_F2A_R_20_13 (.IN_OBUF(tcdm_addr_p2_dup_0[15]),.OUT_OBUF(tcdm_addr_p2[15]));

	qlOBUF QL_INST_F2A_R_20_14 (.IN_OBUF(tcdm_addr_p2_dup_0[16]),.OUT_OBUF(tcdm_addr_p2[16]));

	qlOBUF QL_INST_F2A_R_20_15 (.IN_OBUF(tcdm_addr_p2_dup_0[17]),.OUT_OBUF(tcdm_addr_p2[17]));

	qlOBUF QL_INST_F2A_R_20_16 (.IN_OBUF(tcdm_addr_p2_dup_0[18]),.OUT_OBUF(tcdm_addr_p2[18]));

	qlOBUF QL_INST_F2A_R_20_17 (.IN_OBUF(tcdm_addr_p2_dup_0[19]),.OUT_OBUF(tcdm_addr_p2[19]));

	qlIBUF QL_INST_A2F_R_20_1 (.IN_IBUF(tcdm_rdata_p2[16]),.OUT_IBUF(tcdm_rdata_p2_int[16]));

	qlIBUF QL_INST_A2F_R_20_2 (.IN_IBUF(tcdm_rdata_p2[17]),.OUT_IBUF(tcdm_rdata_p2_int[17]));

	qlIBUF QL_INST_A2F_R_20_3 (.IN_IBUF(tcdm_rdata_p2[18]),.OUT_IBUF(tcdm_rdata_p2_int[18]));

	qlIBUF QL_INST_A2F_R_20_4 (.IN_IBUF(tcdm_rdata_p2[19]),.OUT_IBUF(tcdm_rdata_p2_int[19]));

	qlIBUF QL_INST_A2F_R_20_5 (.IN_IBUF(tcdm_rdata_p2[20]),.OUT_IBUF(tcdm_rdata_p2_int[20]));

	qlIBUF QL_INST_A2F_R_20_6 (.IN_IBUF(tcdm_rdata_p2[21]),.OUT_IBUF(tcdm_rdata_p2_int[21]));

	qlOBUF QL_INST_F2A_R_21_0 (.IN_OBUF(tcdm_wdata_p2_dup_0[24]),.OUT_OBUF(tcdm_wdata_p2[24]));

	qlOBUF QL_INST_F2A_R_21_1 (.IN_OBUF(tcdm_wdata_p2_dup_0[25]),.OUT_OBUF(tcdm_wdata_p2[25]));

	qlOBUF QL_INST_F2A_R_21_2 (.IN_OBUF(tcdm_wdata_p2_dup_0[26]),.OUT_OBUF(tcdm_wdata_p2[26]));

	qlOBUF QL_INST_F2A_R_21_3 (.IN_OBUF(tcdm_wdata_p2_dup_0[27]),.OUT_OBUF(tcdm_wdata_p2[27]));

	qlOBUF QL_INST_F2A_R_21_4 (.IN_OBUF(tcdm_wdata_p2_dup_0[28]),.OUT_OBUF(tcdm_wdata_p2[28]));

	qlOBUF QL_INST_F2A_R_21_5 (.IN_OBUF(tcdm_wdata_p2_dup_0[29]),.OUT_OBUF(tcdm_wdata_p2[29]));

	qlOBUF QL_INST_F2A_R_21_6 (.IN_OBUF(tcdm_wdata_p2_dup_0[30]),.OUT_OBUF(tcdm_wdata_p2[30]));

	qlOBUF QL_INST_F2A_R_21_7 (.IN_OBUF(tcdm_wdata_p2_dup_0[31]),.OUT_OBUF(tcdm_wdata_p2[31]));

	qlIBUF QL_INST_A2F_R_21_0 (.IN_IBUF(tcdm_rdata_p2[22]),.OUT_IBUF(tcdm_rdata_p2_int[22]));

	qlIBUF QL_INST_A2F_R_21_1 (.IN_IBUF(tcdm_rdata_p2[23]),.OUT_IBUF(tcdm_rdata_p2_int[23]));

	qlIBUF QL_INST_A2F_R_21_2 (.IN_IBUF(tcdm_rdata_p2[24]),.OUT_IBUF(tcdm_rdata_p2_int[24]));

	qlIBUF QL_INST_A2F_R_21_3 (.IN_IBUF(tcdm_rdata_p2[25]),.OUT_IBUF(tcdm_rdata_p2_int[25]));

	qlIBUF QL_INST_A2F_R_21_4 (.IN_IBUF(tcdm_rdata_p2[26]),.OUT_IBUF(tcdm_rdata_p2_int[26]));

	qlIBUF QL_INST_A2F_R_21_5 (.IN_IBUF(tcdm_rdata_p2[27]),.OUT_IBUF(tcdm_rdata_p2_int[27]));

	qlIBUF QL_INST_A2F_R_22_0 (.IN_IBUF(tcdm_rdata_p2[28]),.OUT_IBUF(tcdm_rdata_p2_int[28]));

	qlIBUF QL_INST_A2F_R_22_1 (.IN_IBUF(tcdm_rdata_p2[29]),.OUT_IBUF(tcdm_rdata_p2_int[29]));

	qlIBUF QL_INST_A2F_R_22_2 (.IN_IBUF(tcdm_rdata_p2[30]),.OUT_IBUF(tcdm_rdata_p2_int[30]));

	qlIBUF QL_INST_A2F_R_22_3 (.IN_IBUF(tcdm_rdata_p2[31]),.OUT_IBUF(tcdm_rdata_p2_int[31]));

	qlOBUF QL_INST_F2A_R_23_0 (.IN_OBUF(CLK_int_0__CAND0_BRSTR_33_padClk),.OUT_OBUF(tcdm_clk_p3));

	qlOBUF QL_INST_F2A_R_23_1 (.IN_OBUF(tcdm_req_p3_dup_0),.OUT_OBUF(tcdm_req_p3));

	qlOBUF QL_INST_F2A_R_23_2 (.IN_OBUF(tcdm_wen_p3_dup_0),.OUT_OBUF(tcdm_wen_p3));

	qlOBUF QL_INST_F2A_R_23_3 (.IN_OBUF(tcdm_be_p3_dup_0[0]),.OUT_OBUF(tcdm_be_p3[0]));

	qlOBUF QL_INST_F2A_R_23_4 (.IN_OBUF(tcdm_be_p3_dup_0[1]),.OUT_OBUF(tcdm_be_p3[1]));

	qlOBUF QL_INST_F2A_R_23_5 (.IN_OBUF(tcdm_be_p3_dup_0[2]),.OUT_OBUF(tcdm_be_p3[2]));

	qlOBUF QL_INST_F2A_R_23_6 (.IN_OBUF(tcdm_be_p3_dup_0[3]),.OUT_OBUF(tcdm_be_p3[3]));

	qlOBUF QL_INST_F2A_R_23_8 (.IN_OBUF(tcdm_addr_p3_dup_0[0]),.OUT_OBUF(tcdm_addr_p3[0]));

	qlOBUF QL_INST_F2A_R_23_9 (.IN_OBUF(tcdm_addr_p3_dup_0[1]),.OUT_OBUF(tcdm_addr_p3[1]));

	qlOBUF QL_INST_F2A_R_23_10 (.IN_OBUF(tcdm_addr_p3_dup_0[2]),.OUT_OBUF(tcdm_addr_p3[2]));

	qlOBUF QL_INST_F2A_R_23_11 (.IN_OBUF(tcdm_addr_p3_dup_0[3]),.OUT_OBUF(tcdm_addr_p3[3]));

	qlIBUF QL_INST_A2F_R_23_0 (.IN_IBUF(tcdm_rdata_p3[0]),.OUT_IBUF(tcdm_rdata_p3_int[0]));

	qlIBUF QL_INST_A2F_R_23_1 (.IN_IBUF(tcdm_rdata_p3[1]),.OUT_IBUF(tcdm_rdata_p3_int[1]));

	qlIBUF QL_INST_A2F_R_23_2 (.IN_IBUF(tcdm_rdata_p3[2]),.OUT_IBUF(tcdm_rdata_p3_int[2]));

	qlIBUF QL_INST_A2F_R_23_3 (.IN_IBUF(tcdm_rdata_p3[3]),.OUT_IBUF(tcdm_rdata_p3_int[3]));

	qlIBUF QL_INST_A2F_R_23_4 (.IN_IBUF(tcdm_valid_p3),.OUT_IBUF(tcdm_valid_p3_int));

	qlIBUF QL_INST_A2F_R_23_5 (.IN_IBUF(tcdm_gnt_p3),.OUT_IBUF(tcdm_gnt_p3_int));

	qlOBUF QL_INST_F2A_R_24_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[0]),.OUT_OBUF(tcdm_wdata_p3[0]));

	qlOBUF QL_INST_F2A_R_24_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[1]),.OUT_OBUF(tcdm_wdata_p3[1]));

	qlOBUF QL_INST_F2A_R_24_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[2]),.OUT_OBUF(tcdm_wdata_p3[2]));

	qlOBUF QL_INST_F2A_R_24_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[3]),.OUT_OBUF(tcdm_wdata_p3[3]));

	qlOBUF QL_INST_F2A_R_24_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[4]),.OUT_OBUF(tcdm_wdata_p3[4]));

	qlOBUF QL_INST_F2A_R_24_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[5]),.OUT_OBUF(tcdm_wdata_p3[5]));

	qlOBUF QL_INST_F2A_R_24_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[6]),.OUT_OBUF(tcdm_wdata_p3[6]));

	qlOBUF QL_INST_F2A_R_24_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[7]),.OUT_OBUF(tcdm_wdata_p3[7]));

	qlOBUF QL_INST_F2A_R_24_9 (.IN_OBUF(tcdm_addr_p3_dup_0[4]),.OUT_OBUF(tcdm_addr_p3[4]));

	qlOBUF QL_INST_F2A_R_24_10 (.IN_OBUF(tcdm_addr_p3_dup_0[5]),.OUT_OBUF(tcdm_addr_p3[5]));

	qlOBUF QL_INST_F2A_R_24_11 (.IN_OBUF(tcdm_addr_p3_dup_0[6]),.OUT_OBUF(tcdm_addr_p3[6]));

	qlOBUF QL_INST_F2A_R_24_12 (.IN_OBUF(tcdm_addr_p3_dup_0[7]),.OUT_OBUF(tcdm_addr_p3[7]));

	qlOBUF QL_INST_F2A_R_24_13 (.IN_OBUF(tcdm_addr_p3_dup_0[8]),.OUT_OBUF(tcdm_addr_p3[8]));

	qlOBUF QL_INST_F2A_R_24_14 (.IN_OBUF(tcdm_addr_p3_dup_0[9]),.OUT_OBUF(tcdm_addr_p3[9]));

	qlIBUF QL_INST_A2F_R_24_0 (.IN_IBUF(tcdm_rdata_p3[4]),.OUT_IBUF(tcdm_rdata_p3_int[4]));

	qlIBUF QL_INST_A2F_R_24_1 (.IN_IBUF(tcdm_rdata_p3[5]),.OUT_IBUF(tcdm_rdata_p3_int[5]));

	qlIBUF QL_INST_A2F_R_24_2 (.IN_IBUF(tcdm_rdata_p3[6]),.OUT_IBUF(tcdm_rdata_p3_int[6]));

	qlIBUF QL_INST_A2F_R_24_3 (.IN_IBUF(tcdm_rdata_p3[7]),.OUT_IBUF(tcdm_rdata_p3_int[7]));

	qlIBUF QL_INST_A2F_R_24_4 (.IN_IBUF(tcdm_rdata_p3[8]),.OUT_IBUF(tcdm_rdata_p3_int[8]));

	qlIBUF QL_INST_A2F_R_24_5 (.IN_IBUF(tcdm_rdata_p3[9]),.OUT_IBUF(tcdm_rdata_p3_int[9]));

	qlIBUF QL_INST_A2F_R_24_6 (.IN_IBUF(tcdm_rdata_p3[10]),.OUT_IBUF(tcdm_rdata_p3_int[10]));

	qlIBUF QL_INST_A2F_R_24_7 (.IN_IBUF(tcdm_rdata_p3[11]),.OUT_IBUF(tcdm_rdata_p3_int[11]));

	qlOBUF QL_INST_F2A_R_25_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[8]),.OUT_OBUF(tcdm_wdata_p3[8]));

	qlOBUF QL_INST_F2A_R_25_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[9]),.OUT_OBUF(tcdm_wdata_p3[9]));

	qlOBUF QL_INST_F2A_R_25_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[10]),.OUT_OBUF(tcdm_wdata_p3[10]));

	qlOBUF QL_INST_F2A_R_25_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[11]),.OUT_OBUF(tcdm_wdata_p3[11]));

	qlOBUF QL_INST_F2A_R_25_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[12]),.OUT_OBUF(tcdm_wdata_p3[12]));

	qlOBUF QL_INST_F2A_R_25_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[13]),.OUT_OBUF(tcdm_wdata_p3[13]));

	qlOBUF QL_INST_F2A_R_25_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[14]),.OUT_OBUF(tcdm_wdata_p3[14]));

	qlOBUF QL_INST_F2A_R_25_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[15]),.OUT_OBUF(tcdm_wdata_p3[15]));

	qlOBUF QL_INST_F2A_R_25_8 (.IN_OBUF(tcdm_addr_p3_dup_0[10]),.OUT_OBUF(tcdm_addr_p3[10]));

	qlOBUF QL_INST_F2A_R_25_9 (.IN_OBUF(tcdm_addr_p3_dup_0[11]),.OUT_OBUF(tcdm_addr_p3[11]));

	qlOBUF QL_INST_F2A_R_25_10 (.IN_OBUF(tcdm_addr_p3_dup_0[12]),.OUT_OBUF(tcdm_addr_p3[12]));

	qlOBUF QL_INST_F2A_R_25_11 (.IN_OBUF(tcdm_addr_p3_dup_0[13]),.OUT_OBUF(tcdm_addr_p3[13]));

	qlIBUF QL_INST_A2F_R_25_0 (.IN_IBUF(tcdm_rdata_p3[12]),.OUT_IBUF(tcdm_rdata_p3_int[12]));

	qlIBUF QL_INST_A2F_R_25_1 (.IN_IBUF(tcdm_rdata_p3[13]),.OUT_IBUF(tcdm_rdata_p3_int[13]));

	qlIBUF QL_INST_A2F_R_25_2 (.IN_IBUF(tcdm_rdata_p3[14]),.OUT_IBUF(tcdm_rdata_p3_int[14]));

	qlIBUF QL_INST_A2F_R_25_3 (.IN_IBUF(tcdm_rdata_p3[15]),.OUT_IBUF(tcdm_rdata_p3_int[15]));

	qlIBUF QL_INST_A2F_R_25_4 (.IN_IBUF(tcdm_fmo_p3),.OUT_IBUF(tcdm_fmo_p3_int));

	qlOBUF QL_INST_F2A_R_26_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[16]),.OUT_OBUF(tcdm_wdata_p3[16]));

	qlOBUF QL_INST_F2A_R_26_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[17]),.OUT_OBUF(tcdm_wdata_p3[17]));

	qlOBUF QL_INST_F2A_R_26_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[18]),.OUT_OBUF(tcdm_wdata_p3[18]));

	qlOBUF QL_INST_F2A_R_26_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[19]),.OUT_OBUF(tcdm_wdata_p3[19]));

	qlOBUF QL_INST_F2A_R_26_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[20]),.OUT_OBUF(tcdm_wdata_p3[20]));

	qlOBUF QL_INST_F2A_R_26_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[21]),.OUT_OBUF(tcdm_wdata_p3[21]));

	qlOBUF QL_INST_F2A_R_26_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[22]),.OUT_OBUF(tcdm_wdata_p3[22]));

	qlOBUF QL_INST_F2A_R_26_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[23]),.OUT_OBUF(tcdm_wdata_p3[23]));

	qlOBUF QL_INST_F2A_R_26_12 (.IN_OBUF(tcdm_addr_p3_dup_0[14]),.OUT_OBUF(tcdm_addr_p3[14]));

	qlOBUF QL_INST_F2A_R_26_13 (.IN_OBUF(tcdm_addr_p3_dup_0[15]),.OUT_OBUF(tcdm_addr_p3[15]));

	qlOBUF QL_INST_F2A_R_26_14 (.IN_OBUF(tcdm_addr_p3_dup_0[16]),.OUT_OBUF(tcdm_addr_p3[16]));

	qlOBUF QL_INST_F2A_R_26_15 (.IN_OBUF(tcdm_addr_p3_dup_0[17]),.OUT_OBUF(tcdm_addr_p3[17]));

	qlOBUF QL_INST_F2A_R_26_16 (.IN_OBUF(tcdm_addr_p3_dup_0[18]),.OUT_OBUF(tcdm_addr_p3[18]));

	qlOBUF QL_INST_F2A_R_26_17 (.IN_OBUF(tcdm_addr_p3_dup_0[19]),.OUT_OBUF(tcdm_addr_p3[19]));

	qlIBUF QL_INST_A2F_R_26_1 (.IN_IBUF(tcdm_rdata_p3[16]),.OUT_IBUF(tcdm_rdata_p3_int[16]));

	qlIBUF QL_INST_A2F_R_26_2 (.IN_IBUF(tcdm_rdata_p3[17]),.OUT_IBUF(tcdm_rdata_p3_int[17]));

	qlIBUF QL_INST_A2F_R_26_3 (.IN_IBUF(tcdm_rdata_p3[18]),.OUT_IBUF(tcdm_rdata_p3_int[18]));

	qlIBUF QL_INST_A2F_R_26_4 (.IN_IBUF(tcdm_rdata_p3[19]),.OUT_IBUF(tcdm_rdata_p3_int[19]));

	qlIBUF QL_INST_A2F_R_26_5 (.IN_IBUF(tcdm_rdata_p3[20]),.OUT_IBUF(tcdm_rdata_p3_int[20]));

	qlIBUF QL_INST_A2F_R_26_6 (.IN_IBUF(tcdm_rdata_p3[21]),.OUT_IBUF(tcdm_rdata_p3_int[21]));

	qlOBUF QL_INST_F2A_R_27_0 (.IN_OBUF(tcdm_wdata_p3_dup_0[24]),.OUT_OBUF(tcdm_wdata_p3[24]));

	qlOBUF QL_INST_F2A_R_27_1 (.IN_OBUF(tcdm_wdata_p3_dup_0[25]),.OUT_OBUF(tcdm_wdata_p3[25]));

	qlOBUF QL_INST_F2A_R_27_2 (.IN_OBUF(tcdm_wdata_p3_dup_0[26]),.OUT_OBUF(tcdm_wdata_p3[26]));

	qlOBUF QL_INST_F2A_R_27_3 (.IN_OBUF(tcdm_wdata_p3_dup_0[27]),.OUT_OBUF(tcdm_wdata_p3[27]));

	qlOBUF QL_INST_F2A_R_27_4 (.IN_OBUF(tcdm_wdata_p3_dup_0[28]),.OUT_OBUF(tcdm_wdata_p3[28]));

	qlOBUF QL_INST_F2A_R_27_5 (.IN_OBUF(tcdm_wdata_p3_dup_0[29]),.OUT_OBUF(tcdm_wdata_p3[29]));

	qlOBUF QL_INST_F2A_R_27_6 (.IN_OBUF(tcdm_wdata_p3_dup_0[30]),.OUT_OBUF(tcdm_wdata_p3[30]));

	qlOBUF QL_INST_F2A_R_27_7 (.IN_OBUF(tcdm_wdata_p3_dup_0[31]),.OUT_OBUF(tcdm_wdata_p3[31]));

	qlIBUF QL_INST_A2F_R_27_0 (.IN_IBUF(tcdm_rdata_p3[22]),.OUT_IBUF(tcdm_rdata_p3_int[22]));

	qlIBUF QL_INST_A2F_R_27_1 (.IN_IBUF(tcdm_rdata_p3[23]),.OUT_IBUF(tcdm_rdata_p3_int[23]));

	qlIBUF QL_INST_A2F_R_27_2 (.IN_IBUF(tcdm_rdata_p3[24]),.OUT_IBUF(tcdm_rdata_p3_int[24]));

	qlIBUF QL_INST_A2F_R_27_3 (.IN_IBUF(tcdm_rdata_p3[25]),.OUT_IBUF(tcdm_rdata_p3_int[25]));

	qlIBUF QL_INST_A2F_R_27_4 (.IN_IBUF(tcdm_rdata_p3[26]),.OUT_IBUF(tcdm_rdata_p3_int[26]));

	qlIBUF QL_INST_A2F_R_27_5 (.IN_IBUF(tcdm_rdata_p3[27]),.OUT_IBUF(tcdm_rdata_p3_int[27]));

	qlIBUF QL_INST_A2F_R_28_0 (.IN_IBUF(tcdm_rdata_p3[28]),.OUT_IBUF(tcdm_rdata_p3_int[28]));

	qlIBUF QL_INST_A2F_R_28_1 (.IN_IBUF(tcdm_rdata_p3[29]),.OUT_IBUF(tcdm_rdata_p3_int[29]));

	qlIBUF QL_INST_A2F_R_28_2 (.IN_IBUF(tcdm_rdata_p3[30]),.OUT_IBUF(tcdm_rdata_p3_int[30]));

	qlIBUF QL_INST_A2F_R_28_3 (.IN_IBUF(tcdm_rdata_p3[31]),.OUT_IBUF(tcdm_rdata_p3_int[31]));

	qlIBUF QL_INST_A2F_R_29_2 (.IN_IBUF(RESET[1]),.OUT_IBUF(RESET_int[1]));

	qlOBUF QL_INST_F2A_B_2_0 (.IN_OBUF(CLK_int_0__CAND0_BLSBL_2_padClk),.OUT_OBUF(m1_coef_wclk));

	qlOBUF QL_INST_F2A_B_2_1 (.IN_OBUF(m1_oper0_wmode_dup_0[1]),.OUT_OBUF(m1_oper0_wmode[1]));

	qlOBUF QL_INST_F2A_B_2_2 (.IN_OBUF(m1_oper0_wmode_dup_0[0]),.OUT_OBUF(m1_oper0_wmode[0]));

	qlOBUF QL_INST_F2A_B_2_3 (.IN_OBUF(CLK_int_0__CAND0_BLSBL_2_padClk),.OUT_OBUF(m0_oper1_rclk));

	qlOBUF QL_INST_F2A_B_2_4 (.IN_OBUF(m1_oper0_rmode_dup_0[1]),.OUT_OBUF(m1_oper0_rmode[1]));

	qlOBUF QL_INST_F2A_B_2_5 (.IN_OBUF(m1_oper0_rmode_dup_0[0]),.OUT_OBUF(m1_oper0_rmode[0]));

	qlOBUF QL_INST_F2A_B_2_6 (.IN_OBUF(m1_oper0_wdata_dup_0[31]),.OUT_OBUF(m1_oper0_wdata[31]));

	qlOBUF QL_INST_F2A_B_2_7 (.IN_OBUF(m1_oper0_wdata_dup_0[30]),.OUT_OBUF(m1_oper0_wdata[30]));

	qlOBUF QL_INST_F2A_B_2_8 (.IN_OBUF(m1_oper0_wdata_dup_0[29]),.OUT_OBUF(m1_oper0_wdata[29]));

	qlOBUF QL_INST_F2A_B_2_9 (.IN_OBUF(m1_oper0_wdata_dup_0[28]),.OUT_OBUF(m1_oper0_wdata[28]));

	qlOBUF QL_INST_F2A_B_2_10 (.IN_OBUF(m1_oper0_wdata_dup_0[27]),.OUT_OBUF(m1_oper0_wdata[27]));

	qlOBUF QL_INST_F2A_B_2_11 (.IN_OBUF(m1_oper0_wdata_dup_0[26]),.OUT_OBUF(m1_oper0_wdata[26]));

	qlOBUF QL_INST_F2A_B_2_12 (.IN_OBUF(m1_oper0_wdata_dup_0[25]),.OUT_OBUF(m1_oper0_wdata[25]));

	qlOBUF QL_INST_F2A_B_2_13 (.IN_OBUF(m1_oper0_wdata_dup_0[24]),.OUT_OBUF(m1_oper0_wdata[24]));

	qlOBUF QL_INST_F2A_B_2_14 (.IN_OBUF(m1_oper0_wdata_dup_0[23]),.OUT_OBUF(m1_oper0_wdata[23]));

	qlOBUF QL_INST_F2A_B_2_15 (.IN_OBUF(m1_oper0_wdata_dup_0[22]),.OUT_OBUF(m1_oper0_wdata[22]));

	qlOBUF QL_INST_F2A_B_2_16 (.IN_OBUF(m1_oper0_wdata_dup_0[21]),.OUT_OBUF(m1_oper0_wdata[21]));

	qlOBUF QL_INST_F2A_B_2_17 (.IN_OBUF(m1_oper0_wdata_dup_0[20]),.OUT_OBUF(m1_oper0_wdata[20]));

	qlIBUF QL_INST_A2F_B_2_0 (.IN_IBUF(m1_oper0_rdata[31]),.OUT_IBUF(m1_oper0_rdata_int[31]));

	qlIBUF QL_INST_A2F_B_2_1 (.IN_IBUF(m1_oper0_rdata[30]),.OUT_IBUF(m1_oper0_rdata_int[30]));

	qlIBUF QL_INST_A2F_B_2_2 (.IN_IBUF(m1_oper0_rdata[29]),.OUT_IBUF(m1_oper0_rdata_int[29]));

	qlIBUF QL_INST_A2F_B_2_3 (.IN_IBUF(m1_oper0_rdata[28]),.OUT_IBUF(m1_oper0_rdata_int[28]));

	qlOBUF QL_INST_F2A_B_3_0 (.IN_OBUF(m1_oper0_wdata_dup_0[19]),.OUT_OBUF(m1_oper0_wdata[19]));

	qlOBUF QL_INST_F2A_B_3_1 (.IN_OBUF(m1_oper0_wdata_dup_0[18]),.OUT_OBUF(m1_oper0_wdata[18]));

	qlOBUF QL_INST_F2A_B_3_2 (.IN_OBUF(m1_oper0_wdata_dup_0[17]),.OUT_OBUF(m1_oper0_wdata[17]));

	qlOBUF QL_INST_F2A_B_3_3 (.IN_OBUF(m1_oper0_wdata_dup_0[16]),.OUT_OBUF(m1_oper0_wdata[16]));

	qlOBUF QL_INST_F2A_B_3_4 (.IN_OBUF(m1_oper0_wdata_dup_0[15]),.OUT_OBUF(m1_oper0_wdata[15]));

	qlOBUF QL_INST_F2A_B_3_5 (.IN_OBUF(m1_oper0_wdata_dup_0[14]),.OUT_OBUF(m1_oper0_wdata[14]));

	qlOBUF QL_INST_F2A_B_3_6 (.IN_OBUF(m1_oper0_wdata_dup_0[13]),.OUT_OBUF(m1_oper0_wdata[13]));

	qlOBUF QL_INST_F2A_B_3_7 (.IN_OBUF(m1_oper0_wdata_dup_0[12]),.OUT_OBUF(m1_oper0_wdata[12]));

	qlOBUF QL_INST_F2A_B_3_8 (.IN_OBUF(m1_oper0_wdata_dup_0[11]),.OUT_OBUF(m1_oper0_wdata[11]));

	qlOBUF QL_INST_F2A_B_3_9 (.IN_OBUF(m1_oper0_wdata_dup_0[10]),.OUT_OBUF(m1_oper0_wdata[10]));

	qlOBUF QL_INST_F2A_B_3_10 (.IN_OBUF(m1_oper0_wdata_dup_0[9]),.OUT_OBUF(m1_oper0_wdata[9]));

	qlOBUF QL_INST_F2A_B_3_11 (.IN_OBUF(m1_oper0_wdata_dup_0[8]),.OUT_OBUF(m1_oper0_wdata[8]));

	qlIBUF QL_INST_A2F_B_3_0 (.IN_IBUF(m1_oper0_rdata[27]),.OUT_IBUF(m1_oper0_rdata_int[27]));

	qlIBUF QL_INST_A2F_B_3_1 (.IN_IBUF(m1_oper0_rdata[26]),.OUT_IBUF(m1_oper0_rdata_int[26]));

	qlIBUF QL_INST_A2F_B_3_2 (.IN_IBUF(m1_oper0_rdata[25]),.OUT_IBUF(m1_oper0_rdata_int[25]));

	qlIBUF QL_INST_A2F_B_3_3 (.IN_IBUF(m1_oper0_rdata[24]),.OUT_IBUF(m1_oper0_rdata_int[24]));

	qlIBUF QL_INST_A2F_B_3_4 (.IN_IBUF(m1_oper0_rdata[23]),.OUT_IBUF(m1_oper0_rdata_int[23]));

	qlIBUF QL_INST_A2F_B_3_5 (.IN_IBUF(m1_oper0_rdata[22]),.OUT_IBUF(m1_oper0_rdata_int[22]));

	qlOBUF QL_INST_F2A_B_4_0 (.IN_OBUF(m1_oper0_wdata_dup_0[7]),.OUT_OBUF(m1_oper0_wdata[7]));

	qlOBUF QL_INST_F2A_B_4_1 (.IN_OBUF(m1_oper0_wdata_dup_0[6]),.OUT_OBUF(m1_oper0_wdata[6]));

	qlOBUF QL_INST_F2A_B_4_2 (.IN_OBUF(m1_oper0_wdata_dup_0[5]),.OUT_OBUF(m1_oper0_wdata[5]));

	qlOBUF QL_INST_F2A_B_4_3 (.IN_OBUF(m1_oper0_wdata_dup_0[4]),.OUT_OBUF(m1_oper0_wdata[4]));

	qlOBUF QL_INST_F2A_B_4_4 (.IN_OBUF(m1_oper0_wdata_dup_0[3]),.OUT_OBUF(m1_oper0_wdata[3]));

	qlOBUF QL_INST_F2A_B_4_5 (.IN_OBUF(m1_oper0_wdata_dup_0[2]),.OUT_OBUF(m1_oper0_wdata[2]));

	qlOBUF QL_INST_F2A_B_4_6 (.IN_OBUF(m1_oper0_wdata_dup_0[1]),.OUT_OBUF(m1_oper0_wdata[1]));

	qlOBUF QL_INST_F2A_B_4_7 (.IN_OBUF(m1_oper0_wdata_dup_0[0]),.OUT_OBUF(m1_oper0_wdata[0]));

	qlOBUF QL_INST_F2A_B_4_8 (.IN_OBUF(m1_oper0_waddr_dup_0[11]),.OUT_OBUF(m1_oper0_waddr[11]));

	qlOBUF QL_INST_F2A_B_4_9 (.IN_OBUF(m1_oper0_waddr_dup_0[10]),.OUT_OBUF(m1_oper0_waddr[10]));

	qlOBUF QL_INST_F2A_B_4_10 (.IN_OBUF(m1_oper0_waddr_dup_0[9]),.OUT_OBUF(m1_oper0_waddr[9]));

	qlOBUF QL_INST_F2A_B_4_11 (.IN_OBUF(m1_oper0_waddr_dup_0[8]),.OUT_OBUF(m1_oper0_waddr[8]));

	qlOBUF QL_INST_F2A_B_4_12 (.IN_OBUF(m1_oper0_waddr_dup_0[7]),.OUT_OBUF(m1_oper0_waddr[7]));

	qlOBUF QL_INST_F2A_B_4_13 (.IN_OBUF(m1_oper0_waddr_dup_0[6]),.OUT_OBUF(m1_oper0_waddr[6]));

	qlOBUF QL_INST_F2A_B_4_14 (.IN_OBUF(m1_oper0_waddr_dup_0[5]),.OUT_OBUF(m1_oper0_waddr[5]));

	qlOBUF QL_INST_F2A_B_4_15 (.IN_OBUF(m1_oper0_waddr_dup_0[4]),.OUT_OBUF(m1_oper0_waddr[4]));

	qlOBUF QL_INST_F2A_B_4_16 (.IN_OBUF(m1_oper0_waddr_dup_0[3]),.OUT_OBUF(m1_oper0_waddr[3]));

	qlOBUF QL_INST_F2A_B_4_17 (.IN_OBUF(m1_oper0_waddr_dup_0[2]),.OUT_OBUF(m1_oper0_waddr[2]));

	qlIBUF QL_INST_A2F_B_4_0 (.IN_IBUF(m1_oper0_rdata[21]),.OUT_IBUF(m1_oper0_rdata_int[21]));

	qlIBUF QL_INST_A2F_B_4_1 (.IN_IBUF(m1_oper0_rdata[20]),.OUT_IBUF(m1_oper0_rdata_int[20]));

	qlIBUF QL_INST_A2F_B_4_2 (.IN_IBUF(m1_oper0_rdata[19]),.OUT_IBUF(m1_oper0_rdata_int[19]));

	qlIBUF QL_INST_A2F_B_4_3 (.IN_IBUF(m1_oper0_rdata[18]),.OUT_IBUF(m1_oper0_rdata_int[18]));

	qlIBUF QL_INST_A2F_B_4_4 (.IN_IBUF(m1_oper0_rdata[17]),.OUT_IBUF(m1_oper0_rdata_int[17]));

	qlIBUF QL_INST_A2F_B_4_5 (.IN_IBUF(m1_oper0_rdata[16]),.OUT_IBUF(m1_oper0_rdata_int[16]));

	qlIBUF QL_INST_A2F_B_4_6 (.IN_IBUF(m1_oper0_rdata[15]),.OUT_IBUF(m1_oper0_rdata_int[15]));

	qlIBUF QL_INST_A2F_B_4_7 (.IN_IBUF(m1_oper0_rdata[14]),.OUT_IBUF(m1_oper0_rdata_int[14]));

	qlOBUF QL_INST_F2A_B_5_0 (.IN_OBUF(m1_oper0_waddr_dup_0[1]),.OUT_OBUF(m1_oper0_waddr[1]));

	qlOBUF QL_INST_F2A_B_5_1 (.IN_OBUF(m1_oper0_waddr_dup_0[0]),.OUT_OBUF(m1_oper0_waddr[0]));

	qlOBUF QL_INST_F2A_B_5_2 (.IN_OBUF(m0_oper0_wdsel_dup_0),.OUT_OBUF(m0_oper0_wdsel));

	qlOBUF QL_INST_F2A_B_5_3 (.IN_OBUF(m1_oper0_raddr_dup_0[11]),.OUT_OBUF(m1_oper0_raddr[11]));

	qlOBUF QL_INST_F2A_B_5_4 (.IN_OBUF(m1_oper0_raddr_dup_0[10]),.OUT_OBUF(m1_oper0_raddr[10]));

	qlOBUF QL_INST_F2A_B_5_5 (.IN_OBUF(m1_oper0_raddr_dup_0[9]),.OUT_OBUF(m1_oper0_raddr[9]));

	qlOBUF QL_INST_F2A_B_5_6 (.IN_OBUF(m1_oper0_raddr_dup_0[8]),.OUT_OBUF(m1_oper0_raddr[8]));

	qlOBUF QL_INST_F2A_B_5_7 (.IN_OBUF(m1_oper0_raddr_dup_0[7]),.OUT_OBUF(m1_oper0_raddr[7]));

	qlOBUF QL_INST_F2A_B_5_8 (.IN_OBUF(m1_oper0_raddr_dup_0[6]),.OUT_OBUF(m1_oper0_raddr[6]));

	qlOBUF QL_INST_F2A_B_5_9 (.IN_OBUF(m1_oper0_raddr_dup_0[5]),.OUT_OBUF(m1_oper0_raddr[5]));

	qlOBUF QL_INST_F2A_B_5_10 (.IN_OBUF(m1_oper0_raddr_dup_0[4]),.OUT_OBUF(m1_oper0_raddr[4]));

	qlOBUF QL_INST_F2A_B_5_11 (.IN_OBUF(m1_oper0_raddr_dup_0[3]),.OUT_OBUF(m1_oper0_raddr[3]));

	qlIBUF QL_INST_A2F_B_5_0 (.IN_IBUF(m1_oper0_rdata[13]),.OUT_IBUF(m1_oper0_rdata_int[13]));

	qlIBUF QL_INST_A2F_B_5_1 (.IN_IBUF(m1_oper0_rdata[12]),.OUT_IBUF(m1_oper0_rdata_int[12]));

	qlIBUF QL_INST_A2F_B_5_2 (.IN_IBUF(m1_oper0_rdata[11]),.OUT_IBUF(m1_oper0_rdata_int[11]));

	qlIBUF QL_INST_A2F_B_5_3 (.IN_IBUF(m1_oper0_rdata[10]),.OUT_IBUF(m1_oper0_rdata_int[10]));

	qlIBUF QL_INST_A2F_B_5_4 (.IN_IBUF(m1_oper0_rdata[9]),.OUT_IBUF(m1_oper0_rdata_int[9]));

	qlIBUF QL_INST_A2F_B_5_5 (.IN_IBUF(m1_oper0_rdata[8]),.OUT_IBUF(m1_oper0_rdata_int[8]));

	qlOBUF QL_INST_F2A_B_6_0 (.IN_OBUF(m0_m1_sat_dup_0),.OUT_OBUF(m0_m1_sat));

	qlOBUF QL_INST_F2A_B_6_1 (.IN_OBUF(m1_oper0_raddr_dup_0[2]),.OUT_OBUF(m1_oper0_raddr[2]));

	qlOBUF QL_INST_F2A_B_6_2 (.IN_OBUF(GND),.OUT_OBUF(m1_oper0_raddr[1]));

	qlOBUF QL_INST_F2A_B_6_3 (.IN_OBUF(GND),.OUT_OBUF(m1_oper0_raddr[0]));

	qlOBUF QL_INST_F2A_B_6_4 (.IN_OBUF(m1_oper0_we_dup_0),.OUT_OBUF(m1_oper0_we));

	qlOBUF QL_INST_F2A_B_6_5 (.IN_OBUF(m1_m1_clr_dup_0),.OUT_OBUF(m1_m1_clr));

	qlOBUF QL_INST_F2A_B_6_6 (.IN_OBUF(m1_m0_outsel_dup_0[5]),.OUT_OBUF(m1_m0_outsel[5]));

	qlOBUF QL_INST_F2A_B_6_7 (.IN_OBUF(m1_m0_outsel_dup_0[4]),.OUT_OBUF(m1_m0_outsel[4]));

	qlOBUF QL_INST_F2A_B_6_8 (.IN_OBUF(m1_m0_outsel_dup_0[3]),.OUT_OBUF(m1_m0_outsel[3]));

	qlOBUF QL_INST_F2A_B_6_9 (.IN_OBUF(m1_m0_outsel_dup_0[2]),.OUT_OBUF(m1_m0_outsel[2]));

	qlOBUF QL_INST_F2A_B_6_10 (.IN_OBUF(m1_m0_outsel_dup_0[1]),.OUT_OBUF(m1_m0_outsel[1]));

	qlOBUF QL_INST_F2A_B_6_11 (.IN_OBUF(m1_m0_outsel_dup_0[0]),.OUT_OBUF(m1_m0_outsel[0]));

	qlOBUF QL_INST_F2A_B_6_12 (.IN_OBUF(m0_m0_tc_dup_0),.OUT_OBUF(m0_m0_tc));

	qlOBUF QL_INST_F2A_B_6_13 (.IN_OBUF(m0_m0_osel_dup_0),.OUT_OBUF(m0_m0_osel));

	qlOBUF QL_INST_F2A_B_6_14 (.IN_OBUF(m1_m0_tc_dup_0),.OUT_OBUF(m1_m0_tc));

	qlOBUF QL_INST_F2A_B_6_15 (.IN_OBUF(m1_oper0_rdata_int[31]),.OUT_OBUF(m1_m0_oper_in[31]));

	qlOBUF QL_INST_F2A_B_6_16 (.IN_OBUF(m1_oper0_rdata_int[30]),.OUT_OBUF(m1_m0_oper_in[30]));

	qlOBUF QL_INST_F2A_B_6_17 (.IN_OBUF(m1_oper0_rdata_int[29]),.OUT_OBUF(m1_m0_oper_in[29]));

	DBUF QL_INST_F2Adef_B_6_1 (.IN_DBUF(GND),.OUT_DBUF(m1_coef_powerdn));

	qlIBUF QL_INST_A2F_B_6_0 (.IN_IBUF(m1_oper0_rdata[7]),.OUT_IBUF(m1_oper0_rdata_int[7]));

	qlIBUF QL_INST_A2F_B_6_1 (.IN_IBUF(m1_oper0_rdata[6]),.OUT_IBUF(m1_oper0_rdata_int[6]));

	qlIBUF QL_INST_A2F_B_6_2 (.IN_IBUF(m1_oper0_rdata[5]),.OUT_IBUF(m1_oper0_rdata_int[5]));

	qlIBUF QL_INST_A2F_B_6_3 (.IN_IBUF(m1_oper0_rdata[4]),.OUT_IBUF(m1_oper0_rdata_int[4]));

	qlIBUF QL_INST_A2F_B_6_4 (.IN_IBUF(m1_oper0_rdata[3]),.OUT_IBUF(m1_oper0_rdata_int[3]));

	qlIBUF QL_INST_A2F_B_6_5 (.IN_IBUF(m1_oper0_rdata[2]),.OUT_IBUF(m1_oper0_rdata_int[2]));

	qlIBUF QL_INST_A2F_B_6_6 (.IN_IBUF(m1_oper0_rdata[1]),.OUT_IBUF(m1_oper0_rdata_int[1]));

	qlIBUF QL_INST_A2F_B_6_7 (.IN_IBUF(m1_oper0_rdata[0]),.OUT_IBUF(m1_oper0_rdata_int[0]));

	qlOBUF QL_INST_F2A_B_7_0 (.IN_OBUF(m0_m0_csel_dup_0),.OUT_OBUF(m0_m0_csel));

	qlOBUF QL_INST_F2A_B_7_1 (.IN_OBUF(m1_oper0_rdata_int[28]),.OUT_OBUF(m1_m0_oper_in[28]));

	qlOBUF QL_INST_F2A_B_7_2 (.IN_OBUF(m1_oper0_rdata_int[27]),.OUT_OBUF(m1_m0_oper_in[27]));

	qlOBUF QL_INST_F2A_B_7_3 (.IN_OBUF(m1_oper0_rdata_int[26]),.OUT_OBUF(m1_m0_oper_in[26]));

	qlOBUF QL_INST_F2A_B_7_4 (.IN_OBUF(m1_oper0_rdata_int[25]),.OUT_OBUF(m1_m0_oper_in[25]));

	qlOBUF QL_INST_F2A_B_7_5 (.IN_OBUF(m1_oper0_rdata_int[24]),.OUT_OBUF(m1_m0_oper_in[24]));

	qlOBUF QL_INST_F2A_B_7_6 (.IN_OBUF(m1_oper0_rdata_int[23]),.OUT_OBUF(m1_m0_oper_in[23]));

	qlOBUF QL_INST_F2A_B_7_7 (.IN_OBUF(m1_oper0_rdata_int[22]),.OUT_OBUF(m1_m0_oper_in[22]));

	qlOBUF QL_INST_F2A_B_7_8 (.IN_OBUF(m1_oper0_rdata_int[21]),.OUT_OBUF(m1_m0_oper_in[21]));

	qlOBUF QL_INST_F2A_B_7_9 (.IN_OBUF(m1_oper0_rdata_int[20]),.OUT_OBUF(m1_m0_oper_in[20]));

	qlOBUF QL_INST_F2A_B_7_10 (.IN_OBUF(m1_oper0_rdata_int[19]),.OUT_OBUF(m1_m0_oper_in[19]));

	qlOBUF QL_INST_F2A_B_7_11 (.IN_OBUF(m1_oper0_rdata_int[18]),.OUT_OBUF(m1_m0_oper_in[18]));

	qlIBUF QL_INST_A2F_B_7_0 (.IN_IBUF(m1_m0_dataout[31]),.OUT_IBUF(m1_m0_dataout_int[31]));

	qlIBUF QL_INST_A2F_B_7_1 (.IN_IBUF(m1_m0_dataout[30]),.OUT_IBUF(m1_m0_dataout_int[30]));

	qlIBUF QL_INST_A2F_B_7_2 (.IN_IBUF(m1_m0_dataout[29]),.OUT_IBUF(m1_m0_dataout_int[29]));

	qlIBUF QL_INST_A2F_B_7_3 (.IN_IBUF(m1_m0_dataout[28]),.OUT_IBUF(m1_m0_dataout_int[28]));

	qlIBUF QL_INST_A2F_B_7_4 (.IN_IBUF(m1_m0_dataout[27]),.OUT_IBUF(m1_m0_dataout_int[27]));

	qlIBUF QL_INST_A2F_B_7_5 (.IN_IBUF(m1_m0_dataout[26]),.OUT_IBUF(m1_m0_dataout_int[26]));

	qlOBUF QL_INST_F2A_B_8_0 (.IN_OBUF(m1_oper0_rdata_int[17]),.OUT_OBUF(m1_m0_oper_in[17]));

	qlOBUF QL_INST_F2A_B_8_1 (.IN_OBUF(m1_oper0_rdata_int[16]),.OUT_OBUF(m1_m0_oper_in[16]));

	qlOBUF QL_INST_F2A_B_8_2 (.IN_OBUF(m1_oper0_rdata_int[15]),.OUT_OBUF(m1_m0_oper_in[15]));

	qlOBUF QL_INST_F2A_B_8_3 (.IN_OBUF(m1_oper0_rdata_int[14]),.OUT_OBUF(m1_m0_oper_in[14]));

	qlOBUF QL_INST_F2A_B_8_4 (.IN_OBUF(m1_oper0_rdata_int[13]),.OUT_OBUF(m1_m0_oper_in[13]));

	qlOBUF QL_INST_F2A_B_8_5 (.IN_OBUF(m1_oper0_rdata_int[12]),.OUT_OBUF(m1_m0_oper_in[12]));

	qlOBUF QL_INST_F2A_B_8_6 (.IN_OBUF(m1_oper0_rdata_int[11]),.OUT_OBUF(m1_m0_oper_in[11]));

	qlOBUF QL_INST_F2A_B_8_7 (.IN_OBUF(m1_oper0_rdata_int[10]),.OUT_OBUF(m1_m0_oper_in[10]));

	qlOBUF QL_INST_F2A_B_8_8 (.IN_OBUF(m1_oper0_rdata_int[9]),.OUT_OBUF(m1_m0_oper_in[9]));

	qlOBUF QL_INST_F2A_B_8_9 (.IN_OBUF(m1_oper0_rdata_int[8]),.OUT_OBUF(m1_m0_oper_in[8]));

	qlOBUF QL_INST_F2A_B_8_10 (.IN_OBUF(m1_oper0_rdata_int[7]),.OUT_OBUF(m1_m0_oper_in[7]));

	qlOBUF QL_INST_F2A_B_8_11 (.IN_OBUF(m1_oper0_rdata_int[6]),.OUT_OBUF(m1_m0_oper_in[6]));

	qlOBUF QL_INST_F2A_B_8_12 (.IN_OBUF(m1_oper0_rdata_int[5]),.OUT_OBUF(m1_m0_oper_in[5]));

	qlOBUF QL_INST_F2A_B_8_13 (.IN_OBUF(m1_oper0_rdata_int[4]),.OUT_OBUF(m1_m0_oper_in[4]));

	qlOBUF QL_INST_F2A_B_8_14 (.IN_OBUF(m1_oper0_rdata_int[3]),.OUT_OBUF(m1_m0_oper_in[3]));

	qlOBUF QL_INST_F2A_B_8_15 (.IN_OBUF(m1_oper0_rdata_int[2]),.OUT_OBUF(m1_m0_oper_in[2]));

	qlOBUF QL_INST_F2A_B_8_16 (.IN_OBUF(m1_oper0_rdata_int[1]),.OUT_OBUF(m1_m0_oper_in[1]));

	qlOBUF QL_INST_F2A_B_8_17 (.IN_OBUF(m1_oper0_rdata_int[0]),.OUT_OBUF(m1_m0_oper_in[0]));

	qlIBUF QL_INST_A2F_B_8_0 (.IN_IBUF(m1_m0_dataout[25]),.OUT_IBUF(m1_m0_dataout_int[25]));

	qlIBUF QL_INST_A2F_B_8_1 (.IN_IBUF(m1_m0_dataout[24]),.OUT_IBUF(m1_m0_dataout_int[24]));

	qlIBUF QL_INST_A2F_B_8_2 (.IN_IBUF(m1_m0_dataout[23]),.OUT_IBUF(m1_m0_dataout_int[23]));

	qlIBUF QL_INST_A2F_B_8_3 (.IN_IBUF(m1_m0_dataout[22]),.OUT_IBUF(m1_m0_dataout_int[22]));

	qlIBUF QL_INST_A2F_B_8_4 (.IN_IBUF(m1_m0_dataout[21]),.OUT_IBUF(m1_m0_dataout_int[21]));

	qlIBUF QL_INST_A2F_B_8_5 (.IN_IBUF(m1_m0_dataout[20]),.OUT_IBUF(m1_m0_dataout_int[20]));

	qlIBUF QL_INST_A2F_B_8_6 (.IN_IBUF(m1_m0_dataout[19]),.OUT_IBUF(m1_m0_dataout_int[19]));

	qlIBUF QL_INST_A2F_B_8_7 (.IN_IBUF(m1_m0_dataout[18]),.OUT_IBUF(m1_m0_dataout_int[18]));

	qlOBUF QL_INST_F2A_B_9_0 (.IN_OBUF(m1_m1_tc_dup_0),.OUT_OBUF(m1_m1_tc));

	qlOBUF QL_INST_F2A_B_9_1 (.IN_OBUF(m1_coef_rdata_int[31]),.OUT_OBUF(m1_m0_coef_in[31]));

	qlOBUF QL_INST_F2A_B_9_2 (.IN_OBUF(m1_coef_rdata_int[30]),.OUT_OBUF(m1_m0_coef_in[30]));

	qlOBUF QL_INST_F2A_B_9_3 (.IN_OBUF(m1_coef_rdata_int[29]),.OUT_OBUF(m1_m0_coef_in[29]));

	qlOBUF QL_INST_F2A_B_9_4 (.IN_OBUF(m1_coef_rdata_int[28]),.OUT_OBUF(m1_m0_coef_in[28]));

	qlOBUF QL_INST_F2A_B_9_5 (.IN_OBUF(m1_coef_rdata_int[27]),.OUT_OBUF(m1_m0_coef_in[27]));

	qlOBUF QL_INST_F2A_B_9_6 (.IN_OBUF(m1_coef_rdata_int[26]),.OUT_OBUF(m1_m0_coef_in[26]));

	qlOBUF QL_INST_F2A_B_9_7 (.IN_OBUF(m1_coef_rdata_int[25]),.OUT_OBUF(m1_m0_coef_in[25]));

	qlOBUF QL_INST_F2A_B_9_8 (.IN_OBUF(m1_coef_rdata_int[24]),.OUT_OBUF(m1_m0_coef_in[24]));

	qlOBUF QL_INST_F2A_B_9_9 (.IN_OBUF(m1_coef_rdata_int[23]),.OUT_OBUF(m1_m0_coef_in[23]));

	qlOBUF QL_INST_F2A_B_9_10 (.IN_OBUF(m1_coef_rdata_int[22]),.OUT_OBUF(m1_m0_coef_in[22]));

	qlOBUF QL_INST_F2A_B_9_11 (.IN_OBUF(m1_coef_rdata_int[21]),.OUT_OBUF(m1_m0_coef_in[21]));

	qlIBUF QL_INST_A2F_B_9_0 (.IN_IBUF(m1_m0_dataout[17]),.OUT_IBUF(m1_m0_dataout_int[17]));

	qlIBUF QL_INST_A2F_B_9_1 (.IN_IBUF(m1_m0_dataout[16]),.OUT_IBUF(m1_m0_dataout_int[16]));

	qlIBUF QL_INST_A2F_B_9_2 (.IN_IBUF(m1_m0_dataout[15]),.OUT_IBUF(m1_m0_dataout_int[15]));

	qlIBUF QL_INST_A2F_B_9_3 (.IN_IBUF(m1_m0_dataout[14]),.OUT_IBUF(m1_m0_dataout_int[14]));

	qlIBUF QL_INST_A2F_B_9_4 (.IN_IBUF(m1_m0_dataout[13]),.OUT_IBUF(m1_m0_dataout_int[13]));

	qlIBUF QL_INST_A2F_B_9_5 (.IN_IBUF(m1_m0_dataout[12]),.OUT_IBUF(m1_m0_dataout_int[12]));

	qlOBUF QL_INST_F2A_B_10_0 (.IN_OBUF(m1_coef_rdata_int[20]),.OUT_OBUF(m1_m0_coef_in[20]));

	qlOBUF QL_INST_F2A_B_10_1 (.IN_OBUF(m1_coef_rdata_int[19]),.OUT_OBUF(m1_m0_coef_in[19]));

	qlOBUF QL_INST_F2A_B_10_2 (.IN_OBUF(m1_coef_rdata_int[18]),.OUT_OBUF(m1_m0_coef_in[18]));

	qlOBUF QL_INST_F2A_B_10_3 (.IN_OBUF(m1_coef_rdata_int[17]),.OUT_OBUF(m1_m0_coef_in[17]));

	qlOBUF QL_INST_F2A_B_10_4 (.IN_OBUF(m1_coef_rdata_int[16]),.OUT_OBUF(m1_m0_coef_in[16]));

	qlOBUF QL_INST_F2A_B_10_5 (.IN_OBUF(m1_coef_rdata_int[15]),.OUT_OBUF(m1_m0_coef_in[15]));

	qlOBUF QL_INST_F2A_B_10_6 (.IN_OBUF(m1_coef_rdata_int[14]),.OUT_OBUF(m1_m0_coef_in[14]));

	qlOBUF QL_INST_F2A_B_10_7 (.IN_OBUF(m1_coef_rdata_int[13]),.OUT_OBUF(m1_m0_coef_in[13]));

	qlOBUF QL_INST_F2A_B_10_8 (.IN_OBUF(m1_coef_rdata_int[12]),.OUT_OBUF(m1_m0_coef_in[12]));

	qlOBUF QL_INST_F2A_B_10_9 (.IN_OBUF(m1_coef_rdata_int[11]),.OUT_OBUF(m1_m0_coef_in[11]));

	qlOBUF QL_INST_F2A_B_10_10 (.IN_OBUF(m1_coef_rdata_int[10]),.OUT_OBUF(m1_m0_coef_in[10]));

	qlOBUF QL_INST_F2A_B_10_11 (.IN_OBUF(m1_coef_rdata_int[9]),.OUT_OBUF(m1_m0_coef_in[9]));

	qlOBUF QL_INST_F2A_B_10_12 (.IN_OBUF(m1_coef_rdata_int[8]),.OUT_OBUF(m1_m0_coef_in[8]));

	qlOBUF QL_INST_F2A_B_10_13 (.IN_OBUF(m1_coef_rdata_int[7]),.OUT_OBUF(m1_m0_coef_in[7]));

	qlOBUF QL_INST_F2A_B_10_14 (.IN_OBUF(m1_coef_rdata_int[6]),.OUT_OBUF(m1_m0_coef_in[6]));

	qlOBUF QL_INST_F2A_B_10_15 (.IN_OBUF(m1_coef_rdata_int[5]),.OUT_OBUF(m1_m0_coef_in[5]));

	qlOBUF QL_INST_F2A_B_10_16 (.IN_OBUF(m1_coef_rdata_int[4]),.OUT_OBUF(m1_m0_coef_in[4]));

	qlOBUF QL_INST_F2A_B_10_17 (.IN_OBUF(m1_coef_rdata_int[3]),.OUT_OBUF(m1_m0_coef_in[3]));

	qlIBUF QL_INST_A2F_B_10_0 (.IN_IBUF(m1_m0_dataout[11]),.OUT_IBUF(m1_m0_dataout_int[11]));

	qlIBUF QL_INST_A2F_B_10_1 (.IN_IBUF(m1_m0_dataout[10]),.OUT_IBUF(m1_m0_dataout_int[10]));

	qlIBUF QL_INST_A2F_B_10_2 (.IN_IBUF(m1_m0_dataout[9]),.OUT_IBUF(m1_m0_dataout_int[9]));

	qlIBUF QL_INST_A2F_B_10_3 (.IN_IBUF(m1_m0_dataout[8]),.OUT_IBUF(m1_m0_dataout_int[8]));

	qlIBUF QL_INST_A2F_B_10_4 (.IN_IBUF(m1_m0_dataout[7]),.OUT_IBUF(m1_m0_dataout_int[7]));

	qlIBUF QL_INST_A2F_B_10_5 (.IN_IBUF(m1_m0_dataout[6]),.OUT_IBUF(m1_m0_dataout_int[6]));

	qlIBUF QL_INST_A2F_B_10_6 (.IN_IBUF(m1_m0_dataout[5]),.OUT_IBUF(m1_m0_dataout_int[5]));

	qlIBUF QL_INST_A2F_B_10_7 (.IN_IBUF(m1_m0_dataout[4]),.OUT_IBUF(m1_m0_dataout_int[4]));

	qlOBUF QL_INST_F2A_B_11_0 (.IN_OBUF(m1_coef_rdata_int[2]),.OUT_OBUF(m1_m0_coef_in[2]));

	qlOBUF QL_INST_F2A_B_11_1 (.IN_OBUF(m1_coef_rdata_int[1]),.OUT_OBUF(m1_m0_coef_in[1]));

	qlOBUF QL_INST_F2A_B_11_2 (.IN_OBUF(m1_coef_rdata_int[0]),.OUT_OBUF(m1_m0_coef_in[0]));

	qlOBUF QL_INST_F2A_B_11_3 (.IN_OBUF(m1_m0_mode_dup_0[1]),.OUT_OBUF(m1_m0_mode[1]));

	qlOBUF QL_INST_F2A_B_11_4 (.IN_OBUF(m1_m0_mode_dup_0[0]),.OUT_OBUF(m1_m0_mode[0]));

	qlOBUF QL_INST_F2A_B_11_5 (.IN_OBUF(m1_coef_rmode_dup_0[1]),.OUT_OBUF(m1_coef_rmode[1]));

	qlOBUF QL_INST_F2A_B_11_6 (.IN_OBUF(m1_coef_rmode_dup_0[0]),.OUT_OBUF(m1_coef_rmode[0]));

	qlOBUF QL_INST_F2A_B_11_7 (.IN_OBUF(m1_coef_wdata_dup_0[31]),.OUT_OBUF(m1_coef_wdata[31]));

	qlOBUF QL_INST_F2A_B_11_8 (.IN_OBUF(m1_coef_wdata_dup_0[30]),.OUT_OBUF(m1_coef_wdata[30]));

	qlOBUF QL_INST_F2A_B_11_9 (.IN_OBUF(m1_coef_wdata_dup_0[29]),.OUT_OBUF(m1_coef_wdata[29]));

	qlOBUF QL_INST_F2A_B_11_10 (.IN_OBUF(m1_coef_wdata_dup_0[28]),.OUT_OBUF(m1_coef_wdata[28]));

	qlOBUF QL_INST_F2A_B_11_11 (.IN_OBUF(m1_coef_wdata_dup_0[27]),.OUT_OBUF(m1_coef_wdata[27]));

	qlIBUF QL_INST_A2F_B_11_0 (.IN_IBUF(m1_m0_dataout[3]),.OUT_IBUF(m1_m0_dataout_int[3]));

	qlIBUF QL_INST_A2F_B_11_1 (.IN_IBUF(m1_m0_dataout[2]),.OUT_IBUF(m1_m0_dataout_int[2]));

	qlIBUF QL_INST_A2F_B_11_2 (.IN_IBUF(m1_m0_dataout[1]),.OUT_IBUF(m1_m0_dataout_int[1]));

	qlIBUF QL_INST_A2F_B_11_3 (.IN_IBUF(m1_m0_dataout[0]),.OUT_IBUF(m1_m0_dataout_int[0]));

	qlIBUF QL_INST_A2F_B_11_4 (.IN_IBUF(m1_coef_rdata[31]),.OUT_IBUF(m1_coef_rdata_int[31]));

	qlIBUF QL_INST_A2F_B_11_5 (.IN_IBUF(m1_coef_rdata[30]),.OUT_IBUF(m1_coef_rdata_int[30]));

	qlOBUF QL_INST_F2A_B_12_0 (.IN_OBUF(m1_coef_wdata_dup_0[26]),.OUT_OBUF(m1_coef_wdata[26]));

	qlOBUF QL_INST_F2A_B_12_1 (.IN_OBUF(m1_coef_wdata_dup_0[25]),.OUT_OBUF(m1_coef_wdata[25]));

	qlOBUF QL_INST_F2A_B_12_2 (.IN_OBUF(m1_coef_wdata_dup_0[24]),.OUT_OBUF(m1_coef_wdata[24]));

	qlOBUF QL_INST_F2A_B_12_3 (.IN_OBUF(m1_coef_wdata_dup_0[23]),.OUT_OBUF(m1_coef_wdata[23]));

	qlOBUF QL_INST_F2A_B_12_4 (.IN_OBUF(m1_coef_wdata_dup_0[22]),.OUT_OBUF(m1_coef_wdata[22]));

	qlOBUF QL_INST_F2A_B_12_5 (.IN_OBUF(m1_coef_wdata_dup_0[21]),.OUT_OBUF(m1_coef_wdata[21]));

	qlOBUF QL_INST_F2A_B_12_6 (.IN_OBUF(m1_coef_wdata_dup_0[20]),.OUT_OBUF(m1_coef_wdata[20]));

	qlOBUF QL_INST_F2A_B_12_7 (.IN_OBUF(m1_coef_wdata_dup_0[19]),.OUT_OBUF(m1_coef_wdata[19]));

	qlOBUF QL_INST_F2A_B_12_8 (.IN_OBUF(m1_coef_wdata_dup_0[18]),.OUT_OBUF(m1_coef_wdata[18]));

	qlOBUF QL_INST_F2A_B_12_9 (.IN_OBUF(m1_coef_wdata_dup_0[17]),.OUT_OBUF(m1_coef_wdata[17]));

	qlOBUF QL_INST_F2A_B_12_10 (.IN_OBUF(m1_coef_wdata_dup_0[16]),.OUT_OBUF(m1_coef_wdata[16]));

	qlOBUF QL_INST_F2A_B_12_11 (.IN_OBUF(m1_coef_wdata_dup_0[15]),.OUT_OBUF(m1_coef_wdata[15]));

	qlOBUF QL_INST_F2A_B_12_12 (.IN_OBUF(m1_coef_wdata_dup_0[14]),.OUT_OBUF(m1_coef_wdata[14]));

	qlOBUF QL_INST_F2A_B_12_13 (.IN_OBUF(m1_coef_wdata_dup_0[13]),.OUT_OBUF(m1_coef_wdata[13]));

	qlOBUF QL_INST_F2A_B_12_14 (.IN_OBUF(m1_coef_wdata_dup_0[12]),.OUT_OBUF(m1_coef_wdata[12]));

	qlOBUF QL_INST_F2A_B_12_15 (.IN_OBUF(m1_coef_wdata_dup_0[11]),.OUT_OBUF(m1_coef_wdata[11]));

	qlOBUF QL_INST_F2A_B_12_16 (.IN_OBUF(m1_coef_wdata_dup_0[10]),.OUT_OBUF(m1_coef_wdata[10]));

	qlOBUF QL_INST_F2A_B_12_17 (.IN_OBUF(m1_coef_wdata_dup_0[9]),.OUT_OBUF(m1_coef_wdata[9]));

	qlIBUF QL_INST_A2F_B_12_0 (.IN_IBUF(m1_coef_rdata[29]),.OUT_IBUF(m1_coef_rdata_int[29]));

	qlIBUF QL_INST_A2F_B_12_1 (.IN_IBUF(m1_coef_rdata[28]),.OUT_IBUF(m1_coef_rdata_int[28]));

	qlIBUF QL_INST_A2F_B_12_2 (.IN_IBUF(m1_coef_rdata[27]),.OUT_IBUF(m1_coef_rdata_int[27]));

	qlIBUF QL_INST_A2F_B_12_3 (.IN_IBUF(m1_coef_rdata[26]),.OUT_IBUF(m1_coef_rdata_int[26]));

	qlIBUF QL_INST_A2F_B_12_4 (.IN_IBUF(m1_coef_rdata[25]),.OUT_IBUF(m1_coef_rdata_int[25]));

	qlIBUF QL_INST_A2F_B_12_5 (.IN_IBUF(m1_coef_rdata[24]),.OUT_IBUF(m1_coef_rdata_int[24]));

	qlIBUF QL_INST_A2F_B_12_6 (.IN_IBUF(m1_coef_rdata[23]),.OUT_IBUF(m1_coef_rdata_int[23]));

	qlIBUF QL_INST_A2F_B_12_7 (.IN_IBUF(m1_coef_rdata[22]),.OUT_IBUF(m1_coef_rdata_int[22]));

	qlOBUF QL_INST_F2A_B_13_0 (.IN_OBUF(m0_m1_reset_dup_0),.OUT_OBUF(m0_m1_reset));

	qlOBUF QL_INST_F2A_B_13_1 (.IN_OBUF(m1_coef_wdata_dup_0[8]),.OUT_OBUF(m1_coef_wdata[8]));

	qlOBUF QL_INST_F2A_B_13_2 (.IN_OBUF(m1_coef_wdata_dup_0[7]),.OUT_OBUF(m1_coef_wdata[7]));

	qlOBUF QL_INST_F2A_B_13_3 (.IN_OBUF(m1_coef_wdata_dup_0[6]),.OUT_OBUF(m1_coef_wdata[6]));

	qlOBUF QL_INST_F2A_B_13_4 (.IN_OBUF(m1_coef_wdata_dup_0[5]),.OUT_OBUF(m1_coef_wdata[5]));

	qlOBUF QL_INST_F2A_B_13_5 (.IN_OBUF(m1_coef_wdata_dup_0[4]),.OUT_OBUF(m1_coef_wdata[4]));

	qlOBUF QL_INST_F2A_B_13_6 (.IN_OBUF(m1_coef_wdata_dup_0[3]),.OUT_OBUF(m1_coef_wdata[3]));

	qlOBUF QL_INST_F2A_B_13_7 (.IN_OBUF(m1_coef_wdata_dup_0[2]),.OUT_OBUF(m1_coef_wdata[2]));

	qlOBUF QL_INST_F2A_B_13_8 (.IN_OBUF(m1_coef_wdata_dup_0[1]),.OUT_OBUF(m1_coef_wdata[1]));

	qlOBUF QL_INST_F2A_B_13_9 (.IN_OBUF(m1_coef_wdata_dup_0[0]),.OUT_OBUF(m1_coef_wdata[0]));

	qlOBUF QL_INST_F2A_B_13_10 (.IN_OBUF(m1_coef_waddr_dup_0[11]),.OUT_OBUF(m1_coef_waddr[11]));

	qlOBUF QL_INST_F2A_B_13_11 (.IN_OBUF(m1_coef_waddr_dup_0[10]),.OUT_OBUF(m1_coef_waddr[10]));

	DBUF QL_INST_F2Adef_B_13_0 (.IN_DBUF(GND),.OUT_DBUF(m0_coef_powerdn));

	qlIBUF QL_INST_A2F_B_13_0 (.IN_IBUF(m1_coef_rdata[21]),.OUT_IBUF(m1_coef_rdata_int[21]));

	qlIBUF QL_INST_A2F_B_13_1 (.IN_IBUF(m1_coef_rdata[20]),.OUT_IBUF(m1_coef_rdata_int[20]));

	qlIBUF QL_INST_A2F_B_13_2 (.IN_IBUF(m1_coef_rdata[19]),.OUT_IBUF(m1_coef_rdata_int[19]));

	qlIBUF QL_INST_A2F_B_13_3 (.IN_IBUF(m1_coef_rdata[18]),.OUT_IBUF(m1_coef_rdata_int[18]));

	qlIBUF QL_INST_A2F_B_13_4 (.IN_IBUF(m1_coef_rdata[17]),.OUT_IBUF(m1_coef_rdata_int[17]));

	qlIBUF QL_INST_A2F_B_13_5 (.IN_IBUF(m1_coef_rdata[16]),.OUT_IBUF(m1_coef_rdata_int[16]));

	qlOBUF QL_INST_F2A_B_14_0 (.IN_OBUF(m1_coef_waddr_dup_0[9]),.OUT_OBUF(m1_coef_waddr[9]));

	qlOBUF QL_INST_F2A_B_14_1 (.IN_OBUF(m1_coef_waddr_dup_0[8]),.OUT_OBUF(m1_coef_waddr[8]));

	qlOBUF QL_INST_F2A_B_14_2 (.IN_OBUF(m1_coef_waddr_dup_0[7]),.OUT_OBUF(m1_coef_waddr[7]));

	qlOBUF QL_INST_F2A_B_14_3 (.IN_OBUF(m1_coef_waddr_dup_0[6]),.OUT_OBUF(m1_coef_waddr[6]));

	qlOBUF QL_INST_F2A_B_14_4 (.IN_OBUF(m1_coef_waddr_dup_0[5]),.OUT_OBUF(m1_coef_waddr[5]));

	qlOBUF QL_INST_F2A_B_14_5 (.IN_OBUF(m1_coef_waddr_dup_0[4]),.OUT_OBUF(m1_coef_waddr[4]));

	qlOBUF QL_INST_F2A_B_14_6 (.IN_OBUF(m1_coef_waddr_dup_0[3]),.OUT_OBUF(m1_coef_waddr[3]));

	qlOBUF QL_INST_F2A_B_14_7 (.IN_OBUF(m1_coef_waddr_dup_0[2]),.OUT_OBUF(m1_coef_waddr[2]));

	qlOBUF QL_INST_F2A_B_14_8 (.IN_OBUF(m1_coef_waddr_dup_0[1]),.OUT_OBUF(m1_coef_waddr[1]));

	qlOBUF QL_INST_F2A_B_14_9 (.IN_OBUF(m1_coef_waddr_dup_0[0]),.OUT_OBUF(m1_coef_waddr[0]));

	qlOBUF QL_INST_F2A_B_14_10 (.IN_OBUF(m0_coef_wdsel_dup_0),.OUT_OBUF(m0_coef_wdsel));

	qlOBUF QL_INST_F2A_B_14_11 (.IN_OBUF(m1_coef_wdsel_dup_0),.OUT_OBUF(m1_coef_wdsel));

	qlOBUF QL_INST_F2A_B_14_12 (.IN_OBUF(m1_coef_we_dup_0),.OUT_OBUF(m1_coef_we));

	qlOBUF QL_INST_F2A_B_14_13 (.IN_OBUF(m1_m0_clken_dup_0),.OUT_OBUF(m1_m0_clken));

	qlOBUF QL_INST_F2A_B_14_14 (.IN_OBUF(m1_coef_raddr_dup_0[11]),.OUT_OBUF(m1_coef_raddr[11]));

	qlOBUF QL_INST_F2A_B_14_15 (.IN_OBUF(m1_coef_raddr_dup_0[10]),.OUT_OBUF(m1_coef_raddr[10]));

	qlOBUF QL_INST_F2A_B_14_16 (.IN_OBUF(m1_coef_raddr_dup_0[9]),.OUT_OBUF(m1_coef_raddr[9]));

	qlOBUF QL_INST_F2A_B_14_17 (.IN_OBUF(m1_coef_raddr_dup_0[8]),.OUT_OBUF(m1_coef_raddr[8]));

	qlIBUF QL_INST_A2F_B_14_0 (.IN_IBUF(m1_coef_rdata[15]),.OUT_IBUF(m1_coef_rdata_int[15]));

	qlIBUF QL_INST_A2F_B_14_1 (.IN_IBUF(m1_coef_rdata[14]),.OUT_IBUF(m1_coef_rdata_int[14]));

	qlIBUF QL_INST_A2F_B_14_2 (.IN_IBUF(m1_coef_rdata[13]),.OUT_IBUF(m1_coef_rdata_int[13]));

	qlIBUF QL_INST_A2F_B_14_3 (.IN_IBUF(m1_coef_rdata[12]),.OUT_IBUF(m1_coef_rdata_int[12]));

	qlIBUF QL_INST_A2F_B_14_4 (.IN_IBUF(m1_coef_rdata[11]),.OUT_IBUF(m1_coef_rdata_int[11]));

	qlIBUF QL_INST_A2F_B_14_5 (.IN_IBUF(m1_coef_rdata[10]),.OUT_IBUF(m1_coef_rdata_int[10]));

	qlIBUF QL_INST_A2F_B_14_6 (.IN_IBUF(m1_coef_rdata[9]),.OUT_IBUF(m1_coef_rdata_int[9]));

	qlIBUF QL_INST_A2F_B_14_7 (.IN_IBUF(m1_coef_rdata[8]),.OUT_IBUF(m1_coef_rdata_int[8]));

	qlOBUF QL_INST_F2A_B_15_0 (.IN_OBUF(m0_m0_rnd_dup_0),.OUT_OBUF(m0_m0_rnd));

	qlOBUF QL_INST_F2A_B_15_1 (.IN_OBUF(m1_coef_raddr_dup_0[7]),.OUT_OBUF(m1_coef_raddr[7]));

	qlOBUF QL_INST_F2A_B_15_2 (.IN_OBUF(m1_coef_raddr_dup_0[6]),.OUT_OBUF(m1_coef_raddr[6]));

	qlOBUF QL_INST_F2A_B_15_3 (.IN_OBUF(m1_coef_raddr_dup_0[5]),.OUT_OBUF(m1_coef_raddr[5]));

	qlOBUF QL_INST_F2A_B_15_4 (.IN_OBUF(m1_coef_raddr_dup_0[4]),.OUT_OBUF(m1_coef_raddr[4]));

	qlOBUF QL_INST_F2A_B_15_5 (.IN_OBUF(m1_coef_raddr_dup_0[3]),.OUT_OBUF(m1_coef_raddr[3]));

	qlOBUF QL_INST_F2A_B_15_6 (.IN_OBUF(m1_coef_raddr_dup_0[2]),.OUT_OBUF(m1_coef_raddr[2]));

	qlOBUF QL_INST_F2A_B_15_7 (.IN_OBUF(m1_coef_raddr_dup_0[1]),.OUT_OBUF(m1_coef_raddr[1]));

	qlOBUF QL_INST_F2A_B_15_8 (.IN_OBUF(m1_coef_raddr_dup_0[0]),.OUT_OBUF(m1_coef_raddr[0]));

	qlOBUF QL_INST_F2A_B_15_9 (.IN_OBUF(m1_coef_wmode_dup_0[1]),.OUT_OBUF(m1_coef_wmode[1]));

	qlOBUF QL_INST_F2A_B_15_10 (.IN_OBUF(m1_coef_wmode_dup_0[0]),.OUT_OBUF(m1_coef_wmode[0]));

	qlIBUF QL_INST_A2F_B_15_0 (.IN_IBUF(m1_coef_rdata[7]),.OUT_IBUF(m1_coef_rdata_int[7]));

	qlIBUF QL_INST_A2F_B_15_1 (.IN_IBUF(m1_coef_rdata[6]),.OUT_IBUF(m1_coef_rdata_int[6]));

	qlIBUF QL_INST_A2F_B_15_2 (.IN_IBUF(m1_coef_rdata[5]),.OUT_IBUF(m1_coef_rdata_int[5]));

	qlIBUF QL_INST_A2F_B_15_3 (.IN_IBUF(m1_coef_rdata[4]),.OUT_IBUF(m1_coef_rdata_int[4]));

	qlIBUF QL_INST_A2F_B_15_4 (.IN_IBUF(m1_coef_rdata[3]),.OUT_IBUF(m1_coef_rdata_int[3]));

	qlIBUF QL_INST_A2F_B_15_5 (.IN_IBUF(m1_coef_rdata[2]),.OUT_IBUF(m1_coef_rdata_int[2]));

	qlIBUF QL_INST_A2F_B_16_0 (.IN_IBUF(m1_coef_rdata[1]),.OUT_IBUF(m1_coef_rdata_int[1]));

	qlIBUF QL_INST_A2F_B_16_1 (.IN_IBUF(m1_coef_rdata[0]),.OUT_IBUF(m1_coef_rdata_int[0]));

	qlOBUF QL_INST_F2A_B_18_7 (.IN_OBUF(m0_m0_outsel_dup_0[5]),.OUT_OBUF(m1_m1_outsel[5]));

	qlOBUF QL_INST_F2A_B_18_8 (.IN_OBUF(m0_m0_outsel_dup_0[4]),.OUT_OBUF(m1_m1_outsel[4]));

	qlOBUF QL_INST_F2A_B_18_9 (.IN_OBUF(m0_m0_outsel_dup_0[3]),.OUT_OBUF(m1_m1_outsel[3]));

	qlOBUF QL_INST_F2A_B_18_10 (.IN_OBUF(m0_m0_outsel_dup_0[2]),.OUT_OBUF(m1_m1_outsel[2]));

	qlOBUF QL_INST_F2A_B_18_11 (.IN_OBUF(m0_m0_outsel_dup_0[1]),.OUT_OBUF(m1_m1_outsel[1]));

	qlOBUF QL_INST_F2A_B_18_12 (.IN_OBUF(m0_m0_outsel_dup_0[0]),.OUT_OBUF(m1_m1_outsel[0]));

	qlOBUF QL_INST_F2A_B_18_13 (.IN_OBUF(m0_m1_clken_dup_0),.OUT_OBUF(m0_m1_clken));

	qlOBUF QL_INST_F2A_B_18_14 (.IN_OBUF(m0_m0_reset_dup_0),.OUT_OBUF(m0_m0_reset));

	qlOBUF QL_INST_F2A_B_18_15 (.IN_OBUF(m0_m1_osel_dup_0),.OUT_OBUF(m0_m1_osel));

	qlOBUF QL_INST_F2A_B_18_16 (.IN_OBUF(m0_oper1_rmode_dup_0[1]),.OUT_OBUF(m0_oper1_rmode[1]));

	qlIBUF QL_INST_A2F_B_18_6 (.IN_IBUF(m1_m1_dataout[31]),.OUT_IBUF(m1_m1_dataout_int[31]));

	qlIBUF QL_INST_A2F_B_18_7 (.IN_IBUF(m1_m1_dataout[30]),.OUT_IBUF(m1_m1_dataout_int[30]));

	qlOBUF QL_INST_F2A_B_19_0 (.IN_OBUF(m0_oper1_rmode_dup_0[0]),.OUT_OBUF(m0_oper1_rmode[0]));

	qlOBUF QL_INST_F2A_B_19_1 (.IN_OBUF(m0_m1_rnd_dup_0),.OUT_OBUF(m0_m1_rnd));

	qlOBUF QL_INST_F2A_B_19_2 (.IN_OBUF(CLK_int_0__CAND0_BRSBL_19_padClk),.OUT_OBUF(m0_oper1_wclk));

	qlOBUF QL_INST_F2A_B_19_3 (.IN_OBUF(tcdm_wen_p2_dup_0),.OUT_OBUF(tcdm_wen_p2));

	qlOBUF QL_INST_F2A_B_19_4 (.IN_OBUF(m1_coef_rdata_int[31]),.OUT_OBUF(m1_m1_coef_in[31]));

	qlOBUF QL_INST_F2A_B_19_5 (.IN_OBUF(m1_coef_rdata_int[30]),.OUT_OBUF(m1_m1_coef_in[30]));

	qlOBUF QL_INST_F2A_B_19_6 (.IN_OBUF(m1_coef_rdata_int[29]),.OUT_OBUF(m1_m1_coef_in[29]));

	qlOBUF QL_INST_F2A_B_19_7 (.IN_OBUF(m1_coef_rdata_int[28]),.OUT_OBUF(m1_m1_coef_in[28]));

	qlOBUF QL_INST_F2A_B_19_8 (.IN_OBUF(m1_coef_rdata_int[27]),.OUT_OBUF(m1_m1_coef_in[27]));

	qlOBUF QL_INST_F2A_B_19_9 (.IN_OBUF(m1_coef_rdata_int[26]),.OUT_OBUF(m1_m1_coef_in[26]));

	qlOBUF QL_INST_F2A_B_19_10 (.IN_OBUF(m1_coef_rdata_int[25]),.OUT_OBUF(m1_m1_coef_in[25]));

	qlOBUF QL_INST_F2A_B_19_11 (.IN_OBUF(m1_coef_rdata_int[24]),.OUT_OBUF(m1_m1_coef_in[24]));

	qlIBUF QL_INST_A2F_B_19_0 (.IN_IBUF(m1_m1_dataout[29]),.OUT_IBUF(m1_m1_dataout_int[29]));

	qlIBUF QL_INST_A2F_B_19_1 (.IN_IBUF(m1_m1_dataout[28]),.OUT_IBUF(m1_m1_dataout_int[28]));

	qlIBUF QL_INST_A2F_B_19_2 (.IN_IBUF(m1_m1_dataout[27]),.OUT_IBUF(m1_m1_dataout_int[27]));

	qlIBUF QL_INST_A2F_B_19_3 (.IN_IBUF(m1_m1_dataout[26]),.OUT_IBUF(m1_m1_dataout_int[26]));

	qlIBUF QL_INST_A2F_B_19_4 (.IN_IBUF(m1_m1_dataout[25]),.OUT_IBUF(m1_m1_dataout_int[25]));

	qlIBUF QL_INST_A2F_B_19_5 (.IN_IBUF(m1_m1_dataout[24]),.OUT_IBUF(m1_m1_dataout_int[24]));

	qlOBUF QL_INST_F2A_B_20_0 (.IN_OBUF(m1_coef_rdata_int[23]),.OUT_OBUF(m1_m1_coef_in[23]));

	qlOBUF QL_INST_F2A_B_20_1 (.IN_OBUF(m1_coef_rdata_int[22]),.OUT_OBUF(m1_m1_coef_in[22]));

	qlOBUF QL_INST_F2A_B_20_2 (.IN_OBUF(m1_coef_rdata_int[21]),.OUT_OBUF(m1_m1_coef_in[21]));

	qlOBUF QL_INST_F2A_B_20_3 (.IN_OBUF(m1_coef_rdata_int[20]),.OUT_OBUF(m1_m1_coef_in[20]));

	qlOBUF QL_INST_F2A_B_20_4 (.IN_OBUF(m1_coef_rdata_int[19]),.OUT_OBUF(m1_m1_coef_in[19]));

	qlOBUF QL_INST_F2A_B_20_5 (.IN_OBUF(m1_coef_rdata_int[18]),.OUT_OBUF(m1_m1_coef_in[18]));

	qlOBUF QL_INST_F2A_B_20_6 (.IN_OBUF(m1_coef_rdata_int[17]),.OUT_OBUF(m1_m1_coef_in[17]));

	qlOBUF QL_INST_F2A_B_20_7 (.IN_OBUF(m1_coef_rdata_int[16]),.OUT_OBUF(m1_m1_coef_in[16]));

	qlOBUF QL_INST_F2A_B_20_8 (.IN_OBUF(m1_coef_rdata_int[15]),.OUT_OBUF(m1_m1_coef_in[15]));

	qlOBUF QL_INST_F2A_B_20_9 (.IN_OBUF(m1_coef_rdata_int[14]),.OUT_OBUF(m1_m1_coef_in[14]));

	qlOBUF QL_INST_F2A_B_20_10 (.IN_OBUF(m1_coef_rdata_int[13]),.OUT_OBUF(m1_m1_coef_in[13]));

	qlOBUF QL_INST_F2A_B_20_11 (.IN_OBUF(m1_coef_rdata_int[12]),.OUT_OBUF(m1_m1_coef_in[12]));

	qlOBUF QL_INST_F2A_B_20_12 (.IN_OBUF(m1_coef_rdata_int[11]),.OUT_OBUF(m1_m1_coef_in[11]));

	qlOBUF QL_INST_F2A_B_20_13 (.IN_OBUF(m1_coef_rdata_int[10]),.OUT_OBUF(m1_m1_coef_in[10]));

	qlOBUF QL_INST_F2A_B_20_14 (.IN_OBUF(m1_coef_rdata_int[9]),.OUT_OBUF(m1_m1_coef_in[9]));

	qlOBUF QL_INST_F2A_B_20_15 (.IN_OBUF(m1_coef_rdata_int[8]),.OUT_OBUF(m1_m1_coef_in[8]));

	qlOBUF QL_INST_F2A_B_20_16 (.IN_OBUF(m1_coef_rdata_int[7]),.OUT_OBUF(m1_m1_coef_in[7]));

	qlOBUF QL_INST_F2A_B_20_17 (.IN_OBUF(m1_coef_rdata_int[6]),.OUT_OBUF(m1_m1_coef_in[6]));

	qlIBUF QL_INST_A2F_B_20_0 (.IN_IBUF(m1_m1_dataout[23]),.OUT_IBUF(m1_m1_dataout_int[23]));

	qlIBUF QL_INST_A2F_B_20_1 (.IN_IBUF(m1_m1_dataout[22]),.OUT_IBUF(m1_m1_dataout_int[22]));

	qlIBUF QL_INST_A2F_B_20_2 (.IN_IBUF(m1_m1_dataout[21]),.OUT_IBUF(m1_m1_dataout_int[21]));

	qlIBUF QL_INST_A2F_B_20_3 (.IN_IBUF(m1_m1_dataout[20]),.OUT_IBUF(m1_m1_dataout_int[20]));

	qlIBUF QL_INST_A2F_B_20_4 (.IN_IBUF(m1_m1_dataout[19]),.OUT_IBUF(m1_m1_dataout_int[19]));

	qlIBUF QL_INST_A2F_B_20_5 (.IN_IBUF(m1_m1_dataout[18]),.OUT_IBUF(m1_m1_dataout_int[18]));

	qlIBUF QL_INST_A2F_B_20_6 (.IN_IBUF(m1_m1_dataout[17]),.OUT_IBUF(m1_m1_dataout_int[17]));

	qlOBUF QL_INST_F2A_B_21_0 (.IN_OBUF(m1_coef_rdata_int[5]),.OUT_OBUF(m1_m1_coef_in[5]));

	qlOBUF QL_INST_F2A_B_21_1 (.IN_OBUF(m1_coef_rdata_int[4]),.OUT_OBUF(m1_m1_coef_in[4]));

	qlOBUF QL_INST_F2A_B_21_2 (.IN_OBUF(m1_coef_rdata_int[3]),.OUT_OBUF(m1_m1_coef_in[3]));

	qlOBUF QL_INST_F2A_B_21_3 (.IN_OBUF(m1_coef_rdata_int[2]),.OUT_OBUF(m1_m1_coef_in[2]));

	qlOBUF QL_INST_F2A_B_21_4 (.IN_OBUF(m1_coef_rdata_int[1]),.OUT_OBUF(m1_m1_coef_in[1]));

	qlOBUF QL_INST_F2A_B_21_5 (.IN_OBUF(m1_coef_rdata_int[0]),.OUT_OBUF(m1_m1_coef_in[0]));

	qlOBUF QL_INST_F2A_B_21_6 (.IN_OBUF(m1_m1_mode_dup_0[1]),.OUT_OBUF(m1_m1_mode[1]));

	qlOBUF QL_INST_F2A_B_21_7 (.IN_OBUF(m1_oper1_we_dup_0),.OUT_OBUF(m1_oper1_we));

	qlOBUF QL_INST_F2A_B_21_8 (.IN_OBUF(m1_m1_mode_dup_0[0]),.OUT_OBUF(m1_m1_mode[0]));

	qlOBUF QL_INST_F2A_B_21_9 (.IN_OBUF(m1_oper1_rdata_int[31]),.OUT_OBUF(m1_m1_oper_in[31]));

	qlOBUF QL_INST_F2A_B_21_10 (.IN_OBUF(m1_oper1_rdata_int[30]),.OUT_OBUF(m1_m1_oper_in[30]));

	qlOBUF QL_INST_F2A_B_21_11 (.IN_OBUF(m1_oper1_rdata_int[29]),.OUT_OBUF(m1_m1_oper_in[29]));

	qlIBUF QL_INST_A2F_B_21_0 (.IN_IBUF(m1_m1_dataout[16]),.OUT_IBUF(m1_m1_dataout_int[16]));

	qlIBUF QL_INST_A2F_B_21_1 (.IN_IBUF(m1_m1_dataout[15]),.OUT_IBUF(m1_m1_dataout_int[15]));

	qlIBUF QL_INST_A2F_B_21_2 (.IN_IBUF(m1_m1_dataout[14]),.OUT_IBUF(m1_m1_dataout_int[14]));

	qlIBUF QL_INST_A2F_B_21_3 (.IN_IBUF(m1_m1_dataout[13]),.OUT_IBUF(m1_m1_dataout_int[13]));

	qlIBUF QL_INST_A2F_B_21_4 (.IN_IBUF(m1_m1_dataout[12]),.OUT_IBUF(m1_m1_dataout_int[12]));

	qlIBUF QL_INST_A2F_B_21_5 (.IN_IBUF(m1_m1_dataout[11]),.OUT_IBUF(m1_m1_dataout_int[11]));

	qlOBUF QL_INST_F2A_B_22_0 (.IN_OBUF(m1_oper1_rdata_int[28]),.OUT_OBUF(m1_m1_oper_in[28]));

	qlOBUF QL_INST_F2A_B_22_1 (.IN_OBUF(m1_oper1_rdata_int[27]),.OUT_OBUF(m1_m1_oper_in[27]));

	qlOBUF QL_INST_F2A_B_22_2 (.IN_OBUF(m1_oper1_rdata_int[26]),.OUT_OBUF(m1_m1_oper_in[26]));

	qlOBUF QL_INST_F2A_B_22_3 (.IN_OBUF(m1_oper1_rdata_int[25]),.OUT_OBUF(m1_m1_oper_in[25]));

	qlOBUF QL_INST_F2A_B_22_4 (.IN_OBUF(m1_oper1_rdata_int[24]),.OUT_OBUF(m1_m1_oper_in[24]));

	qlOBUF QL_INST_F2A_B_22_5 (.IN_OBUF(m1_oper1_rdata_int[23]),.OUT_OBUF(m1_m1_oper_in[23]));

	qlOBUF QL_INST_F2A_B_22_6 (.IN_OBUF(m1_oper1_rdata_int[22]),.OUT_OBUF(m1_m1_oper_in[22]));

	qlOBUF QL_INST_F2A_B_22_7 (.IN_OBUF(m1_oper1_rdata_int[21]),.OUT_OBUF(m1_m1_oper_in[21]));

	qlOBUF QL_INST_F2A_B_22_8 (.IN_OBUF(m1_oper1_rdata_int[20]),.OUT_OBUF(m1_m1_oper_in[20]));

	qlOBUF QL_INST_F2A_B_22_9 (.IN_OBUF(m1_oper1_rdata_int[19]),.OUT_OBUF(m1_m1_oper_in[19]));

	qlOBUF QL_INST_F2A_B_22_10 (.IN_OBUF(m1_oper1_rdata_int[18]),.OUT_OBUF(m1_m1_oper_in[18]));

	qlOBUF QL_INST_F2A_B_22_11 (.IN_OBUF(m1_oper1_rdata_int[17]),.OUT_OBUF(m1_m1_oper_in[17]));

	qlOBUF QL_INST_F2A_B_22_12 (.IN_OBUF(m1_oper1_rdata_int[16]),.OUT_OBUF(m1_m1_oper_in[16]));

	qlOBUF QL_INST_F2A_B_22_13 (.IN_OBUF(m1_oper1_rdata_int[15]),.OUT_OBUF(m1_m1_oper_in[15]));

	qlOBUF QL_INST_F2A_B_22_14 (.IN_OBUF(m1_oper1_rdata_int[14]),.OUT_OBUF(m1_m1_oper_in[14]));

	qlOBUF QL_INST_F2A_B_22_15 (.IN_OBUF(m1_oper1_rdata_int[13]),.OUT_OBUF(m1_m1_oper_in[13]));

	qlOBUF QL_INST_F2A_B_22_16 (.IN_OBUF(m1_oper1_rdata_int[12]),.OUT_OBUF(m1_m1_oper_in[12]));

	qlOBUF QL_INST_F2A_B_22_17 (.IN_OBUF(m1_oper1_rdata_int[11]),.OUT_OBUF(m1_m1_oper_in[11]));

	qlIBUF QL_INST_A2F_B_22_0 (.IN_IBUF(m1_m1_dataout[10]),.OUT_IBUF(m1_m1_dataout_int[10]));

	qlIBUF QL_INST_A2F_B_22_1 (.IN_IBUF(m1_m1_dataout[9]),.OUT_IBUF(m1_m1_dataout_int[9]));

	qlIBUF QL_INST_A2F_B_22_2 (.IN_IBUF(m1_m1_dataout[8]),.OUT_IBUF(m1_m1_dataout_int[8]));

	qlIBUF QL_INST_A2F_B_22_3 (.IN_IBUF(m1_m1_dataout[7]),.OUT_IBUF(m1_m1_dataout_int[7]));

	qlIBUF QL_INST_A2F_B_22_4 (.IN_IBUF(m1_m1_dataout[6]),.OUT_IBUF(m1_m1_dataout_int[6]));

	qlIBUF QL_INST_A2F_B_22_5 (.IN_IBUF(m1_m1_dataout[5]),.OUT_IBUF(m1_m1_dataout_int[5]));

	qlOBUF QL_INST_F2A_B_23_0 (.IN_OBUF(m1_oper1_rdata_int[10]),.OUT_OBUF(m1_m1_oper_in[10]));

	qlOBUF QL_INST_F2A_B_23_1 (.IN_OBUF(m1_oper1_rdata_int[9]),.OUT_OBUF(m1_m1_oper_in[9]));

	qlOBUF QL_INST_F2A_B_23_2 (.IN_OBUF(m1_oper1_rdata_int[8]),.OUT_OBUF(m1_m1_oper_in[8]));

	qlOBUF QL_INST_F2A_B_23_3 (.IN_OBUF(m1_oper1_rdata_int[7]),.OUT_OBUF(m1_m1_oper_in[7]));

	qlOBUF QL_INST_F2A_B_23_4 (.IN_OBUF(m1_oper1_rdata_int[6]),.OUT_OBUF(m1_m1_oper_in[6]));

	qlOBUF QL_INST_F2A_B_23_5 (.IN_OBUF(m1_oper1_rdata_int[5]),.OUT_OBUF(m1_m1_oper_in[5]));

	qlOBUF QL_INST_F2A_B_23_6 (.IN_OBUF(m1_oper1_rdata_int[4]),.OUT_OBUF(m1_m1_oper_in[4]));

	qlOBUF QL_INST_F2A_B_23_7 (.IN_OBUF(m1_oper1_rdata_int[3]),.OUT_OBUF(m1_m1_oper_in[3]));

	qlOBUF QL_INST_F2A_B_23_8 (.IN_OBUF(m1_oper1_rdata_int[2]),.OUT_OBUF(m1_m1_oper_in[2]));

	qlOBUF QL_INST_F2A_B_23_9 (.IN_OBUF(m1_oper1_rdata_int[1]),.OUT_OBUF(m1_m1_oper_in[1]));

	qlOBUF QL_INST_F2A_B_23_10 (.IN_OBUF(m1_oper1_rdata_int[0]),.OUT_OBUF(m1_m1_oper_in[0]));

	qlIBUF QL_INST_A2F_B_23_0 (.IN_IBUF(m1_m1_dataout[4]),.OUT_IBUF(m1_m1_dataout_int[4]));

	qlIBUF QL_INST_A2F_B_23_1 (.IN_IBUF(m1_m1_dataout[3]),.OUT_IBUF(m1_m1_dataout_int[3]));

	qlIBUF QL_INST_A2F_B_23_2 (.IN_IBUF(m1_m1_dataout[2]),.OUT_IBUF(m1_m1_dataout_int[2]));

	qlIBUF QL_INST_A2F_B_23_3 (.IN_IBUF(m1_m1_dataout[1]),.OUT_IBUF(m1_m1_dataout_int[1]));

	qlIBUF QL_INST_A2F_B_23_4 (.IN_IBUF(m1_m1_dataout[0]),.OUT_IBUF(m1_m1_dataout_int[0]));

	qlOBUF QL_INST_F2A_B_24_16 (.IN_OBUF(m1_oper1_wdata_dup_0[31]),.OUT_OBUF(m1_oper1_wdata[31]));

	qlOBUF QL_INST_F2A_B_24_17 (.IN_OBUF(m1_oper1_wdata_dup_0[30]),.OUT_OBUF(m1_oper1_wdata[30]));

	DBUF QL_INST_F2Adef_B_24_1 (.IN_DBUF(GND),.OUT_DBUF(m0_oper0_powerdn));

	qlOBUF QL_INST_F2A_B_25_0 (.IN_OBUF(m1_oper1_wdata_dup_0[29]),.OUT_OBUF(m1_oper1_wdata[29]));

	qlOBUF QL_INST_F2A_B_25_1 (.IN_OBUF(m1_oper1_wdata_dup_0[28]),.OUT_OBUF(m1_oper1_wdata[28]));

	qlOBUF QL_INST_F2A_B_25_2 (.IN_OBUF(m1_oper1_wdata_dup_0[27]),.OUT_OBUF(m1_oper1_wdata[27]));

	qlOBUF QL_INST_F2A_B_25_3 (.IN_OBUF(m1_oper1_wdata_dup_0[26]),.OUT_OBUF(m1_oper1_wdata[26]));

	qlOBUF QL_INST_F2A_B_25_4 (.IN_OBUF(m1_oper1_wdata_dup_0[25]),.OUT_OBUF(m1_oper1_wdata[25]));

	qlOBUF QL_INST_F2A_B_25_5 (.IN_OBUF(m1_oper1_wdata_dup_0[24]),.OUT_OBUF(m1_oper1_wdata[24]));

	qlOBUF QL_INST_F2A_B_25_6 (.IN_OBUF(m1_oper1_wdata_dup_0[23]),.OUT_OBUF(m1_oper1_wdata[23]));

	qlOBUF QL_INST_F2A_B_25_7 (.IN_OBUF(m1_oper1_wdata_dup_0[22]),.OUT_OBUF(m1_oper1_wdata[22]));

	qlOBUF QL_INST_F2A_B_25_8 (.IN_OBUF(m1_oper1_wdata_dup_0[21]),.OUT_OBUF(m1_oper1_wdata[21]));

	qlOBUF QL_INST_F2A_B_25_9 (.IN_OBUF(m1_oper1_wdata_dup_0[20]),.OUT_OBUF(m1_oper1_wdata[20]));

	qlOBUF QL_INST_F2A_B_25_10 (.IN_OBUF(m1_oper1_wdata_dup_0[19]),.OUT_OBUF(m1_oper1_wdata[19]));

	qlOBUF QL_INST_F2A_B_25_11 (.IN_OBUF(m1_oper1_wdata_dup_0[18]),.OUT_OBUF(m1_oper1_wdata[18]));

	qlIBUF QL_INST_A2F_B_25_1 (.IN_IBUF(m1_oper1_rdata[31]),.OUT_IBUF(m1_oper1_rdata_int[31]));

	qlIBUF QL_INST_A2F_B_25_2 (.IN_IBUF(m1_oper1_rdata[30]),.OUT_IBUF(m1_oper1_rdata_int[30]));

	qlIBUF QL_INST_A2F_B_25_3 (.IN_IBUF(m1_oper1_rdata[29]),.OUT_IBUF(m1_oper1_rdata_int[29]));

	qlIBUF QL_INST_A2F_B_25_4 (.IN_IBUF(m1_oper1_rdata[28]),.OUT_IBUF(m1_oper1_rdata_int[28]));

	qlIBUF QL_INST_A2F_B_25_5 (.IN_IBUF(m1_oper1_rdata[27]),.OUT_IBUF(m1_oper1_rdata_int[27]));

	qlOBUF QL_INST_F2A_B_26_0 (.IN_OBUF(m1_oper1_wdata_dup_0[17]),.OUT_OBUF(m1_oper1_wdata[17]));

	qlOBUF QL_INST_F2A_B_26_1 (.IN_OBUF(m1_oper1_wdata_dup_0[16]),.OUT_OBUF(m1_oper1_wdata[16]));

	qlOBUF QL_INST_F2A_B_26_2 (.IN_OBUF(m1_oper1_wdata_dup_0[15]),.OUT_OBUF(m1_oper1_wdata[15]));

	qlOBUF QL_INST_F2A_B_26_3 (.IN_OBUF(m1_oper1_wdata_dup_0[14]),.OUT_OBUF(m1_oper1_wdata[14]));

	qlOBUF QL_INST_F2A_B_26_4 (.IN_OBUF(m1_oper1_wdata_dup_0[13]),.OUT_OBUF(m1_oper1_wdata[13]));

	qlOBUF QL_INST_F2A_B_26_5 (.IN_OBUF(m1_oper1_wdata_dup_0[12]),.OUT_OBUF(m1_oper1_wdata[12]));

	qlOBUF QL_INST_F2A_B_26_6 (.IN_OBUF(m1_oper1_wdata_dup_0[11]),.OUT_OBUF(m1_oper1_wdata[11]));

	qlOBUF QL_INST_F2A_B_26_7 (.IN_OBUF(m1_oper1_wdata_dup_0[10]),.OUT_OBUF(m1_oper1_wdata[10]));

	qlOBUF QL_INST_F2A_B_26_8 (.IN_OBUF(m1_oper1_wdata_dup_0[9]),.OUT_OBUF(m1_oper1_wdata[9]));

	qlOBUF QL_INST_F2A_B_26_9 (.IN_OBUF(m1_oper1_wdata_dup_0[8]),.OUT_OBUF(m1_oper1_wdata[8]));

	qlOBUF QL_INST_F2A_B_26_10 (.IN_OBUF(m1_oper1_wdata_dup_0[7]),.OUT_OBUF(m1_oper1_wdata[7]));

	qlOBUF QL_INST_F2A_B_26_11 (.IN_OBUF(m1_oper1_wdata_dup_0[6]),.OUT_OBUF(m1_oper1_wdata[6]));

	qlOBUF QL_INST_F2A_B_26_12 (.IN_OBUF(m1_oper1_wdata_dup_0[5]),.OUT_OBUF(m1_oper1_wdata[5]));

	qlOBUF QL_INST_F2A_B_26_13 (.IN_OBUF(m1_oper1_wdata_dup_0[4]),.OUT_OBUF(m1_oper1_wdata[4]));

	qlOBUF QL_INST_F2A_B_26_14 (.IN_OBUF(m1_oper1_wdata_dup_0[3]),.OUT_OBUF(m1_oper1_wdata[3]));

	qlOBUF QL_INST_F2A_B_26_15 (.IN_OBUF(m1_oper1_wdata_dup_0[2]),.OUT_OBUF(m1_oper1_wdata[2]));

	qlOBUF QL_INST_F2A_B_26_16 (.IN_OBUF(m1_oper1_wdata_dup_0[1]),.OUT_OBUF(m1_oper1_wdata[1]));

	qlOBUF QL_INST_F2A_B_26_17 (.IN_OBUF(m1_oper1_wdata_dup_0[0]),.OUT_OBUF(m1_oper1_wdata[0]));

	qlIBUF QL_INST_A2F_B_26_0 (.IN_IBUF(m1_oper1_rdata[26]),.OUT_IBUF(m1_oper1_rdata_int[26]));

	qlIBUF QL_INST_A2F_B_26_1 (.IN_IBUF(m1_oper1_rdata[25]),.OUT_IBUF(m1_oper1_rdata_int[25]));

	qlIBUF QL_INST_A2F_B_26_2 (.IN_IBUF(m1_oper1_rdata[24]),.OUT_IBUF(m1_oper1_rdata_int[24]));

	qlIBUF QL_INST_A2F_B_26_3 (.IN_IBUF(m1_oper1_rdata[23]),.OUT_IBUF(m1_oper1_rdata_int[23]));

	qlIBUF QL_INST_A2F_B_26_4 (.IN_IBUF(m1_oper1_rdata[22]),.OUT_IBUF(m1_oper1_rdata_int[22]));

	qlIBUF QL_INST_A2F_B_26_5 (.IN_IBUF(m1_oper1_rdata[21]),.OUT_IBUF(m1_oper1_rdata_int[21]));

	qlIBUF QL_INST_A2F_B_26_6 (.IN_IBUF(m1_oper1_rdata[20]),.OUT_IBUF(m1_oper1_rdata_int[20]));

	qlIBUF QL_INST_A2F_B_26_7 (.IN_IBUF(m1_oper1_rdata[19]),.OUT_IBUF(m1_oper1_rdata_int[19]));

	qlOBUF QL_INST_F2A_B_27_0 (.IN_OBUF(m1_oper1_waddr_dup_0[11]),.OUT_OBUF(m1_oper1_waddr[11]));

	qlOBUF QL_INST_F2A_B_27_1 (.IN_OBUF(m1_oper1_waddr_dup_0[10]),.OUT_OBUF(m1_oper1_waddr[10]));

	qlOBUF QL_INST_F2A_B_27_2 (.IN_OBUF(m1_oper1_waddr_dup_0[9]),.OUT_OBUF(m1_oper1_waddr[9]));

	qlOBUF QL_INST_F2A_B_27_3 (.IN_OBUF(m1_oper1_waddr_dup_0[8]),.OUT_OBUF(m1_oper1_waddr[8]));

	qlOBUF QL_INST_F2A_B_27_4 (.IN_OBUF(m1_oper1_waddr_dup_0[7]),.OUT_OBUF(m1_oper1_waddr[7]));

	qlOBUF QL_INST_F2A_B_27_5 (.IN_OBUF(m1_oper1_waddr_dup_0[6]),.OUT_OBUF(m1_oper1_waddr[6]));

	qlOBUF QL_INST_F2A_B_27_6 (.IN_OBUF(m1_oper1_waddr_dup_0[5]),.OUT_OBUF(m1_oper1_waddr[5]));

	qlOBUF QL_INST_F2A_B_27_7 (.IN_OBUF(m1_oper1_waddr_dup_0[4]),.OUT_OBUF(m1_oper1_waddr[4]));

	qlOBUF QL_INST_F2A_B_27_8 (.IN_OBUF(m1_oper1_waddr_dup_0[3]),.OUT_OBUF(m1_oper1_waddr[3]));

	qlOBUF QL_INST_F2A_B_27_9 (.IN_OBUF(m1_oper1_waddr_dup_0[2]),.OUT_OBUF(m1_oper1_waddr[2]));

	qlOBUF QL_INST_F2A_B_27_10 (.IN_OBUF(m1_oper1_waddr_dup_0[1]),.OUT_OBUF(m1_oper1_waddr[1]));

	qlOBUF QL_INST_F2A_B_27_11 (.IN_OBUF(m1_oper1_waddr_dup_0[0]),.OUT_OBUF(m1_oper1_waddr[0]));

	qlIBUF QL_INST_A2F_B_27_0 (.IN_IBUF(m1_oper1_rdata[18]),.OUT_IBUF(m1_oper1_rdata_int[18]));

	qlIBUF QL_INST_A2F_B_27_1 (.IN_IBUF(m1_oper1_rdata[17]),.OUT_IBUF(m1_oper1_rdata_int[17]));

	qlIBUF QL_INST_A2F_B_27_2 (.IN_IBUF(m1_oper1_rdata[16]),.OUT_IBUF(m1_oper1_rdata_int[16]));

	qlIBUF QL_INST_A2F_B_27_3 (.IN_IBUF(m1_oper1_rdata[15]),.OUT_IBUF(m1_oper1_rdata_int[15]));

	qlIBUF QL_INST_A2F_B_27_4 (.IN_IBUF(m1_oper1_rdata[14]),.OUT_IBUF(m1_oper1_rdata_int[14]));

	qlIBUF QL_INST_A2F_B_27_5 (.IN_IBUF(m1_oper1_rdata[13]),.OUT_IBUF(m1_oper1_rdata_int[13]));

	qlOBUF QL_INST_F2A_B_28_0 (.IN_OBUF(CLK_int_0__CAND0_BRSBR_28_padClk),.OUT_OBUF(m1_m1_clk));

	qlOBUF QL_INST_F2A_B_28_1 (.IN_OBUF(m1_oper1_wmode_dup_0[1]),.OUT_OBUF(m1_oper1_wmode[1]));

	qlOBUF QL_INST_F2A_B_28_2 (.IN_OBUF(m1_oper1_wmode_dup_0[0]),.OUT_OBUF(m1_oper1_wmode[0]));

	qlOBUF QL_INST_F2A_B_28_4 (.IN_OBUF(CLK_int_0__CAND0_BRSBR_28_padClk),.OUT_OBUF(m1_m0_clk));

	qlOBUF QL_INST_F2A_B_28_15 (.IN_OBUF(m1_oper1_rmode_dup_0[1]),.OUT_OBUF(m1_oper1_rmode[1]));

	qlOBUF QL_INST_F2A_B_28_16 (.IN_OBUF(m1_oper1_rmode_dup_0[0]),.OUT_OBUF(m1_oper1_rmode[0]));

	qlOBUF QL_INST_F2A_B_28_17 (.IN_OBUF(m1_oper1_raddr_dup_0[11]),.OUT_OBUF(m1_oper1_raddr[11]));

	qlIBUF QL_INST_A2F_B_28_1 (.IN_IBUF(m1_oper1_rdata[12]),.OUT_IBUF(m1_oper1_rdata_int[12]));

	qlIBUF QL_INST_A2F_B_28_2 (.IN_IBUF(m1_oper1_rdata[11]),.OUT_IBUF(m1_oper1_rdata_int[11]));

	qlIBUF QL_INST_A2F_B_28_3 (.IN_IBUF(m1_oper1_rdata[10]),.OUT_IBUF(m1_oper1_rdata_int[10]));

	qlIBUF QL_INST_A2F_B_28_4 (.IN_IBUF(m1_oper1_rdata[9]),.OUT_IBUF(m1_oper1_rdata_int[9]));

	qlIBUF QL_INST_A2F_B_28_5 (.IN_IBUF(m1_oper1_rdata[8]),.OUT_IBUF(m1_oper1_rdata_int[8]));

	qlIBUF QL_INST_A2F_B_28_6 (.IN_IBUF(m1_oper1_rdata[7]),.OUT_IBUF(m1_oper1_rdata_int[7]));

	qlIBUF QL_INST_A2F_B_28_7 (.IN_IBUF(m1_oper1_rdata[6]),.OUT_IBUF(m1_oper1_rdata_int[6]));

	qlOBUF QL_INST_F2A_B_29_0 (.IN_OBUF(CLK_int_0__CAND0_BRSBR_29_padClk),.OUT_OBUF(m1_oper0_wclk));

	qlOBUF QL_INST_F2A_B_29_1 (.IN_OBUF(m1_oper1_raddr_dup_0[10]),.OUT_OBUF(m1_oper1_raddr[10]));

	qlOBUF QL_INST_F2A_B_29_2 (.IN_OBUF(m1_oper1_raddr_dup_0[9]),.OUT_OBUF(m1_oper1_raddr[9]));

	qlOBUF QL_INST_F2A_B_29_3 (.IN_OBUF(m1_oper1_raddr_dup_0[8]),.OUT_OBUF(m1_oper1_raddr[8]));

	qlOBUF QL_INST_F2A_B_29_4 (.IN_OBUF(m1_oper1_raddr_dup_0[7]),.OUT_OBUF(m1_oper1_raddr[7]));

	qlOBUF QL_INST_F2A_B_29_5 (.IN_OBUF(m1_oper1_raddr_dup_0[6]),.OUT_OBUF(m1_oper1_raddr[6]));

	qlOBUF QL_INST_F2A_B_29_6 (.IN_OBUF(m1_oper1_raddr_dup_0[5]),.OUT_OBUF(m1_oper1_raddr[5]));

	qlOBUF QL_INST_F2A_B_29_7 (.IN_OBUF(m1_oper1_raddr_dup_0[4]),.OUT_OBUF(m1_oper1_raddr[4]));

	qlOBUF QL_INST_F2A_B_29_8 (.IN_OBUF(m1_oper1_raddr_dup_0[3]),.OUT_OBUF(m1_oper1_raddr[3]));

	qlOBUF QL_INST_F2A_B_29_9 (.IN_OBUF(m1_oper1_raddr_dup_0[2]),.OUT_OBUF(m1_oper1_raddr[2]));

	qlOBUF QL_INST_F2A_B_29_10 (.IN_OBUF(GND),.OUT_OBUF(m1_oper1_raddr[1]));

	qlOBUF QL_INST_F2A_B_29_11 (.IN_OBUF(GND),.OUT_OBUF(m1_oper1_raddr[0]));

	qlIBUF QL_INST_A2F_B_29_0 (.IN_IBUF(m1_oper1_rdata[5]),.OUT_IBUF(m1_oper1_rdata_int[5]));

	qlIBUF QL_INST_A2F_B_29_1 (.IN_IBUF(m1_oper1_rdata[4]),.OUT_IBUF(m1_oper1_rdata_int[4]));

	qlIBUF QL_INST_A2F_B_29_2 (.IN_IBUF(m1_oper1_rdata[3]),.OUT_IBUF(m1_oper1_rdata_int[3]));

	qlIBUF QL_INST_A2F_B_29_3 (.IN_IBUF(m1_oper1_rdata[2]),.OUT_IBUF(m1_oper1_rdata_int[2]));

	qlIBUF QL_INST_A2F_B_29_4 (.IN_IBUF(m1_oper1_rdata[1]),.OUT_IBUF(m1_oper1_rdata_int[1]));

	qlIBUF QL_INST_A2F_B_29_5 (.IN_IBUF(m1_oper1_rdata[0]),.OUT_IBUF(m1_oper1_rdata_int[0]));

	qlOBUF QL_INST_F2A_L_2_0 (.IN_OBUF(fpgaio_out_dup_0[0]),.OUT_OBUF(fpgaio_out[0]));

	qlOBUF QL_INST_F2A_L_2_1 (.IN_OBUF(fpgaio_oe_dup_0[0]),.OUT_OBUF(fpgaio_oe[0]));

	qlOBUF QL_INST_F2A_L_2_2 (.IN_OBUF(fpgaio_out_dup_0[1]),.OUT_OBUF(fpgaio_out[1]));

	qlOBUF QL_INST_F2A_L_2_3 (.IN_OBUF(fpgaio_oe_dup_0[1]),.OUT_OBUF(fpgaio_oe[1]));

	qlOBUF QL_INST_F2A_L_2_4 (.IN_OBUF(fpgaio_out_dup_0[2]),.OUT_OBUF(fpgaio_out[2]));

	qlOBUF QL_INST_F2A_L_2_5 (.IN_OBUF(fpgaio_oe_dup_0[2]),.OUT_OBUF(fpgaio_oe[2]));

	qlOBUF QL_INST_F2A_L_2_6 (.IN_OBUF(fpgaio_out_dup_0[3]),.OUT_OBUF(fpgaio_out[3]));

	qlOBUF QL_INST_F2A_L_2_7 (.IN_OBUF(fpgaio_oe_dup_0[3]),.OUT_OBUF(fpgaio_oe[3]));

	qlOBUF QL_INST_F2A_L_2_8 (.IN_OBUF(fpgaio_in_int[0]),.OUT_OBUF(events_o[0]));

	DBUF QL_INST_F2Adef_L_2_0 (.IN_DBUF(VCC),.OUT_DBUF(version[0]));

	DBUF QL_INST_F2Adef_L_2_1 (.IN_DBUF(GND),.OUT_DBUF(version[1]));

	DBUF QL_INST_F2Adef_L_2_2 (.IN_DBUF(VCC),.OUT_DBUF(version[2]));

	DBUF QL_INST_F2Adef_L_2_3 (.IN_DBUF(GND),.OUT_DBUF(version[3]));

	DBUF QL_INST_F2Adef_L_2_4 (.IN_DBUF(VCC),.OUT_DBUF(version[4]));

	DBUF QL_INST_F2Adef_L_2_5 (.IN_DBUF(GND),.OUT_DBUF(version[5]));

	DBUF QL_INST_F2Adef_L_2_6 (.IN_DBUF(VCC),.OUT_DBUF(version[6]));

	qlIBUF QL_INST_A2F_L_2_0 (.IN_IBUF(fpgaio_in[0]),.OUT_IBUF(fpgaio_in_int[0]));

	qlIBUF QL_INST_A2F_L_2_1 (.IN_IBUF(fpgaio_in[1]),.OUT_IBUF(fpgaio_in_int[1]));

	qlIBUF QL_INST_A2F_L_2_2 (.IN_IBUF(fpgaio_in[2]),.OUT_IBUF(fpgaio_in_int[2]));

	qlIBUF QL_INST_A2F_L_2_3 (.IN_IBUF(fpgaio_in[3]),.OUT_IBUF(fpgaio_in_int[3]));

	qlIBUF QL_INST_A2F_L_2_4 (.IN_IBUF(RESET[3]),.OUT_IBUF(RESET_int[3]));

	qlOBUF QL_INST_F2A_L_3_0 (.IN_OBUF(fpgaio_out_dup_0[4]),.OUT_OBUF(fpgaio_out[4]));

	qlOBUF QL_INST_F2A_L_3_1 (.IN_OBUF(fpgaio_oe_dup_0[4]),.OUT_OBUF(fpgaio_oe[4]));

	qlOBUF QL_INST_F2A_L_3_2 (.IN_OBUF(fpgaio_out_dup_0[5]),.OUT_OBUF(fpgaio_out[5]));

	qlOBUF QL_INST_F2A_L_3_3 (.IN_OBUF(fpgaio_oe_dup_0[5]),.OUT_OBUF(fpgaio_oe[5]));

	qlOBUF QL_INST_F2A_L_3_4 (.IN_OBUF(fpgaio_out_dup_0[6]),.OUT_OBUF(fpgaio_out[6]));

	qlOBUF QL_INST_F2A_L_3_5 (.IN_OBUF(fpgaio_oe_dup_0[6]),.OUT_OBUF(fpgaio_oe[6]));

	qlOBUF QL_INST_F2A_L_3_6 (.IN_OBUF(fpgaio_out_dup_0[7]),.OUT_OBUF(fpgaio_out[7]));

	qlOBUF QL_INST_F2A_L_3_7 (.IN_OBUF(fpgaio_oe_dup_0[7]),.OUT_OBUF(fpgaio_oe[7]));

	qlOBUF QL_INST_F2A_L_3_8 (.IN_OBUF(fpgaio_in_int[1]),.OUT_OBUF(events_o[1]));

	qlIBUF QL_INST_A2F_L_3_0 (.IN_IBUF(fpgaio_in[4]),.OUT_IBUF(fpgaio_in_int[4]));

	qlIBUF QL_INST_A2F_L_3_1 (.IN_IBUF(fpgaio_in[5]),.OUT_IBUF(fpgaio_in_int[5]));

	qlIBUF QL_INST_A2F_L_3_2 (.IN_IBUF(fpgaio_in[6]),.OUT_IBUF(fpgaio_in_int[6]));

	qlIBUF QL_INST_A2F_L_3_3 (.IN_IBUF(fpgaio_in[7]),.OUT_IBUF(fpgaio_in_int[7]));

	qlIBUF QL_INST_A2F_L_3_4 (.IN_IBUF(fpgaio_in[8]),.OUT_IBUF(fpgaio_in_int[8]));

	qlIBUF QL_INST_A2F_L_3_5 (.IN_IBUF(fpgaio_in[9]),.OUT_IBUF(fpgaio_in_int[9]));

	qlOBUF QL_INST_F2A_L_4_0 (.IN_OBUF(fpgaio_out_dup_0[8]),.OUT_OBUF(fpgaio_out[8]));

	qlOBUF QL_INST_F2A_L_4_1 (.IN_OBUF(fpgaio_oe_dup_0[8]),.OUT_OBUF(fpgaio_oe[8]));

	qlOBUF QL_INST_F2A_L_4_2 (.IN_OBUF(fpgaio_out_dup_0[9]),.OUT_OBUF(fpgaio_out[9]));

	qlOBUF QL_INST_F2A_L_4_3 (.IN_OBUF(fpgaio_oe_dup_0[9]),.OUT_OBUF(fpgaio_oe[9]));

	qlOBUF QL_INST_F2A_L_4_4 (.IN_OBUF(fpgaio_out_dup_0[10]),.OUT_OBUF(fpgaio_out[10]));

	qlOBUF QL_INST_F2A_L_4_5 (.IN_OBUF(fpgaio_oe_dup_0[10]),.OUT_OBUF(fpgaio_oe[10]));

	qlOBUF QL_INST_F2A_L_4_6 (.IN_OBUF(fpgaio_out_dup_0[11]),.OUT_OBUF(fpgaio_out[11]));

	qlOBUF QL_INST_F2A_L_4_7 (.IN_OBUF(fpgaio_oe_dup_0[11]),.OUT_OBUF(fpgaio_oe[11]));

	qlOBUF QL_INST_F2A_L_4_8 (.IN_OBUF(fpgaio_in_int[2]),.OUT_OBUF(events_o[2]));

	qlOBUF QL_INST_F2A_L_4_9 (.IN_OBUF(fpgaio_out_dup_0[12]),.OUT_OBUF(fpgaio_out[12]));

	qlOBUF QL_INST_F2A_L_4_10 (.IN_OBUF(fpgaio_oe_dup_0[12]),.OUT_OBUF(fpgaio_oe[12]));

	qlOBUF QL_INST_F2A_L_4_11 (.IN_OBUF(fpgaio_out_dup_0[13]),.OUT_OBUF(fpgaio_out[13]));

	qlOBUF QL_INST_F2A_L_4_12 (.IN_OBUF(fpgaio_oe_dup_0[13]),.OUT_OBUF(fpgaio_oe[13]));

	qlOBUF QL_INST_F2A_L_4_13 (.IN_OBUF(fpgaio_out_dup_0[14]),.OUT_OBUF(fpgaio_out[14]));

	qlOBUF QL_INST_F2A_L_4_14 (.IN_OBUF(fpgaio_oe_dup_0[14]),.OUT_OBUF(fpgaio_oe[14]));

	DBUF QL_INST_F2Adef_L_4_0 (.IN_DBUF(GND),.OUT_DBUF(version[7]));

	qlIBUF QL_INST_A2F_L_4_2 (.IN_IBUF(fpgaio_in[10]),.OUT_IBUF(fpgaio_in_int[10]));

	qlIBUF QL_INST_A2F_L_4_3 (.IN_IBUF(fpgaio_in[11]),.OUT_IBUF(fpgaio_in_int[11]));

	qlIBUF QL_INST_A2F_L_4_4 (.IN_IBUF(fpgaio_in[12]),.OUT_IBUF(fpgaio_in_int[12]));

	qlIBUF QL_INST_A2F_L_4_5 (.IN_IBUF(fpgaio_in[13]),.OUT_IBUF(fpgaio_in_int[13]));

	qlIBUF QL_INST_A2F_L_4_6 (.IN_IBUF(fpgaio_in[14]),.OUT_IBUF(fpgaio_in_int[14]));

	qlIBUF QL_INST_A2F_L_4_7 (.IN_IBUF(fpgaio_in[15]),.OUT_IBUF(fpgaio_in_int[15]));

	qlOBUF QL_INST_F2A_L_5_0 (.IN_OBUF(fpgaio_out_dup_0[15]),.OUT_OBUF(fpgaio_out[15]));

	qlOBUF QL_INST_F2A_L_5_1 (.IN_OBUF(fpgaio_oe_dup_0[15]),.OUT_OBUF(fpgaio_oe[15]));

	qlOBUF QL_INST_F2A_L_5_2 (.IN_OBUF(fpgaio_in_int[3]),.OUT_OBUF(events_o[3]));

	qlOBUF QL_INST_F2A_L_5_3 (.IN_OBUF(fpgaio_out_dup_0[16]),.OUT_OBUF(fpgaio_out[16]));

	qlOBUF QL_INST_F2A_L_5_4 (.IN_OBUF(fpgaio_oe_dup_0[16]),.OUT_OBUF(fpgaio_oe[16]));

	qlOBUF QL_INST_F2A_L_5_5 (.IN_OBUF(fpgaio_out_dup_0[17]),.OUT_OBUF(fpgaio_out[17]));

	qlOBUF QL_INST_F2A_L_5_6 (.IN_OBUF(fpgaio_oe_dup_0[17]),.OUT_OBUF(fpgaio_oe[17]));

	qlOBUF QL_INST_F2A_L_5_7 (.IN_OBUF(fpgaio_out_dup_0[18]),.OUT_OBUF(fpgaio_out[18]));

	qlOBUF QL_INST_F2A_L_5_8 (.IN_OBUF(fpgaio_oe_dup_0[18]),.OUT_OBUF(fpgaio_oe[18]));

	qlOBUF QL_INST_F2A_L_5_9 (.IN_OBUF(fpgaio_out_dup_0[19]),.OUT_OBUF(fpgaio_out[19]));

	qlOBUF QL_INST_F2A_L_5_10 (.IN_OBUF(fpgaio_oe_dup_0[19]),.OUT_OBUF(fpgaio_oe[19]));

	qlOBUF QL_INST_F2A_L_5_11 (.IN_OBUF(fpgaio_in_int[4]),.OUT_OBUF(events_o[4]));

	qlIBUF QL_INST_A2F_L_5_0 (.IN_IBUF(fpgaio_in[16]),.OUT_IBUF(fpgaio_in_int[16]));

	qlIBUF QL_INST_A2F_L_5_1 (.IN_IBUF(fpgaio_in[17]),.OUT_IBUF(fpgaio_in_int[17]));

	qlIBUF QL_INST_A2F_L_5_2 (.IN_IBUF(fpgaio_in[18]),.OUT_IBUF(fpgaio_in_int[18]));

	qlIBUF QL_INST_A2F_L_5_3 (.IN_IBUF(fpgaio_in[19]),.OUT_IBUF(fpgaio_in_int[19]));

	qlIBUF QL_INST_A2F_L_5_4 (.IN_IBUF(fpgaio_in[20]),.OUT_IBUF(fpgaio_in_int[20]));

	qlIBUF QL_INST_A2F_L_5_5 (.IN_IBUF(fpgaio_in[21]),.OUT_IBUF(fpgaio_in_int[21]));

	qlOBUF QL_INST_F2A_L_6_0 (.IN_OBUF(fpgaio_out_dup_0[20]),.OUT_OBUF(fpgaio_out[20]));

	qlOBUF QL_INST_F2A_L_6_1 (.IN_OBUF(fpgaio_oe_dup_0[20]),.OUT_OBUF(fpgaio_oe[20]));

	qlOBUF QL_INST_F2A_L_6_2 (.IN_OBUF(fpgaio_out_dup_0[21]),.OUT_OBUF(fpgaio_out[21]));

	qlOBUF QL_INST_F2A_L_6_3 (.IN_OBUF(fpgaio_oe_dup_0[21]),.OUT_OBUF(fpgaio_oe[21]));

	qlOBUF QL_INST_F2A_L_6_4 (.IN_OBUF(fpgaio_out_dup_0[22]),.OUT_OBUF(fpgaio_out[22]));

	qlOBUF QL_INST_F2A_L_6_5 (.IN_OBUF(fpgaio_oe_dup_0[22]),.OUT_OBUF(fpgaio_oe[22]));

	qlOBUF QL_INST_F2A_L_6_6 (.IN_OBUF(fpgaio_out_dup_0[23]),.OUT_OBUF(fpgaio_out[23]));

	qlOBUF QL_INST_F2A_L_6_7 (.IN_OBUF(fpgaio_oe_dup_0[23]),.OUT_OBUF(fpgaio_oe[23]));

	qlOBUF QL_INST_F2A_L_6_8 (.IN_OBUF(fpgaio_in_int[5]),.OUT_OBUF(events_o[5]));

	qlOBUF QL_INST_F2A_L_6_9 (.IN_OBUF(fpgaio_out_dup_0[24]),.OUT_OBUF(fpgaio_out[24]));

	qlOBUF QL_INST_F2A_L_6_10 (.IN_OBUF(fpgaio_oe_dup_0[24]),.OUT_OBUF(fpgaio_oe[24]));

	qlOBUF QL_INST_F2A_L_6_11 (.IN_OBUF(fpgaio_out_dup_0[25]),.OUT_OBUF(fpgaio_out[25]));

	qlOBUF QL_INST_F2A_L_6_12 (.IN_OBUF(fpgaio_oe_dup_0[25]),.OUT_OBUF(fpgaio_oe[25]));

	qlOBUF QL_INST_F2A_L_6_13 (.IN_OBUF(fpgaio_out_dup_0[26]),.OUT_OBUF(fpgaio_out[26]));

	qlOBUF QL_INST_F2A_L_6_14 (.IN_OBUF(fpgaio_oe_dup_0[26]),.OUT_OBUF(fpgaio_oe[26]));

	qlOBUF QL_INST_F2A_L_6_15 (.IN_OBUF(fpgaio_out_dup_0[27]),.OUT_OBUF(fpgaio_out[27]));

	qlOBUF QL_INST_F2A_L_6_16 (.IN_OBUF(fpgaio_oe_dup_0[27]),.OUT_OBUF(fpgaio_oe[27]));

	qlOBUF QL_INST_F2A_L_6_17 (.IN_OBUF(fpgaio_in_int[6]),.OUT_OBUF(events_o[6]));

	qlIBUF QL_INST_A2F_L_6_0 (.IN_IBUF(fpgaio_in[22]),.OUT_IBUF(fpgaio_in_int[22]));

	qlIBUF QL_INST_A2F_L_6_1 (.IN_IBUF(fpgaio_in[23]),.OUT_IBUF(fpgaio_in_int[23]));

	qlIBUF QL_INST_A2F_L_6_2 (.IN_IBUF(fpgaio_in[24]),.OUT_IBUF(fpgaio_in_int[24]));

	qlIBUF QL_INST_A2F_L_6_3 (.IN_IBUF(fpgaio_in[25]),.OUT_IBUF(fpgaio_in_int[25]));

	qlIBUF QL_INST_A2F_L_6_4 (.IN_IBUF(fpgaio_in[26]),.OUT_IBUF(fpgaio_in_int[26]));

	qlIBUF QL_INST_A2F_L_6_5 (.IN_IBUF(fpgaio_in[27]),.OUT_IBUF(fpgaio_in_int[27]));

	qlIBUF QL_INST_A2F_L_7_0 (.IN_IBUF(fpgaio_in[28]),.OUT_IBUF(fpgaio_in_int[28]));

	qlIBUF QL_INST_A2F_L_7_1 (.IN_IBUF(fpgaio_in[29]),.OUT_IBUF(fpgaio_in_int[29]));

	qlIBUF QL_INST_A2F_L_7_2 (.IN_IBUF(fpgaio_in[30]),.OUT_IBUF(fpgaio_in_int[30]));

	qlIBUF QL_INST_A2F_L_7_3 (.IN_IBUF(fpgaio_in[31]),.OUT_IBUF(fpgaio_in_int[31]));

	qlIBUF QL_INST_A2F_L_7_4 (.IN_IBUF(lint_WDATA[0]),.OUT_IBUF(lint_WDATA_int[0]));

	qlIBUF QL_INST_A2F_L_7_5 (.IN_IBUF(lint_WDATA[1]),.OUT_IBUF(lint_WDATA_int[1]));

	qlOBUF QL_INST_F2A_L_8_0 (.IN_OBUF(fpgaio_out_dup_0[28]),.OUT_OBUF(fpgaio_out[28]));

	qlOBUF QL_INST_F2A_L_8_1 (.IN_OBUF(fpgaio_oe_dup_0[28]),.OUT_OBUF(fpgaio_oe[28]));

	qlOBUF QL_INST_F2A_L_8_2 (.IN_OBUF(fpgaio_out_dup_0[29]),.OUT_OBUF(fpgaio_out[29]));

	qlOBUF QL_INST_F2A_L_8_3 (.IN_OBUF(fpgaio_oe_dup_0[29]),.OUT_OBUF(fpgaio_oe[29]));

	qlOBUF QL_INST_F2A_L_8_4 (.IN_OBUF(fpgaio_out_dup_0[30]),.OUT_OBUF(fpgaio_out[30]));

	qlOBUF QL_INST_F2A_L_8_5 (.IN_OBUF(fpgaio_oe_dup_0[30]),.OUT_OBUF(fpgaio_oe[30]));

	qlOBUF QL_INST_F2A_L_8_6 (.IN_OBUF(fpgaio_out_dup_0[31]),.OUT_OBUF(fpgaio_out[31]));

	qlOBUF QL_INST_F2A_L_8_7 (.IN_OBUF(fpgaio_oe_dup_0[31]),.OUT_OBUF(fpgaio_oe[31]));

	qlOBUF QL_INST_F2A_L_8_8 (.IN_OBUF(fpgaio_in_int[7]),.OUT_OBUF(events_o[7]));

	qlIBUF QL_INST_A2F_L_8_0 (.IN_IBUF(lint_WDATA[2]),.OUT_IBUF(lint_WDATA_int[2]));

	qlIBUF QL_INST_A2F_L_8_1 (.IN_IBUF(lint_WDATA[3]),.OUT_IBUF(lint_WDATA_int[3]));

	qlIBUF QL_INST_A2F_L_8_2 (.IN_IBUF(lint_WDATA[4]),.OUT_IBUF(lint_WDATA_int[4]));

	qlIBUF QL_INST_A2F_L_8_3 (.IN_IBUF(lint_WDATA[5]),.OUT_IBUF(lint_WDATA_int[5]));

	qlIBUF QL_INST_A2F_L_8_4 (.IN_IBUF(lint_WDATA[6]),.OUT_IBUF(lint_WDATA_int[6]));

	qlIBUF QL_INST_A2F_L_8_5 (.IN_IBUF(lint_WDATA[7]),.OUT_IBUF(lint_WDATA_int[7]));

	qlIBUF QL_INST_A2F_L_8_6 (.IN_IBUF(lint_WDATA[8]),.OUT_IBUF(lint_WDATA_int[8]));

	qlIBUF QL_INST_A2F_L_8_7 (.IN_IBUF(lint_WDATA[9]),.OUT_IBUF(lint_WDATA_int[9]));

	qlIBUF QL_INST_A2F_L_9_0 (.IN_IBUF(lint_WDATA[10]),.OUT_IBUF(lint_WDATA_int[10]));

	qlIBUF QL_INST_A2F_L_9_1 (.IN_IBUF(lint_WDATA[11]),.OUT_IBUF(lint_WDATA_int[11]));

	qlIBUF QL_INST_A2F_L_9_2 (.IN_IBUF(lint_WDATA[12]),.OUT_IBUF(lint_WDATA_int[12]));

	qlIBUF QL_INST_A2F_L_9_3 (.IN_IBUF(lint_WDATA[13]),.OUT_IBUF(lint_WDATA_int[13]));

	qlIBUF QL_INST_A2F_L_9_4 (.IN_IBUF(lint_WDATA[14]),.OUT_IBUF(lint_WDATA_int[14]));

	qlIBUF QL_INST_A2F_L_9_5 (.IN_IBUF(lint_WDATA[15]),.OUT_IBUF(lint_WDATA_int[15]));

	qlIBUF QL_INST_A2F_L_10_0 (.IN_IBUF(lint_WDATA[16]),.OUT_IBUF(lint_WDATA_int[16]));

	qlIBUF QL_INST_A2F_L_10_1 (.IN_IBUF(lint_WDATA[17]),.OUT_IBUF(lint_WDATA_int[17]));

	qlIBUF QL_INST_A2F_L_10_2 (.IN_IBUF(lint_WDATA[18]),.OUT_IBUF(lint_WDATA_int[18]));

	qlIBUF QL_INST_A2F_L_10_3 (.IN_IBUF(lint_WDATA[19]),.OUT_IBUF(lint_WDATA_int[19]));

	qlIBUF QL_INST_A2F_L_10_4 (.IN_IBUF(lint_WDATA[20]),.OUT_IBUF(lint_WDATA_int[20]));

	qlIBUF QL_INST_A2F_L_10_5 (.IN_IBUF(lint_WDATA[21]),.OUT_IBUF(lint_WDATA_int[21]));

	qlIBUF QL_INST_A2F_L_10_6 (.IN_IBUF(lint_WDATA[22]),.OUT_IBUF(lint_WDATA_int[22]));

	qlIBUF QL_INST_A2F_L_10_7 (.IN_IBUF(lint_WDATA[23]),.OUT_IBUF(lint_WDATA_int[23]));

	qlIBUF QL_INST_A2F_L_11_0 (.IN_IBUF(lint_WDATA[24]),.OUT_IBUF(lint_WDATA_int[24]));

	qlIBUF QL_INST_A2F_L_11_1 (.IN_IBUF(lint_WDATA[25]),.OUT_IBUF(lint_WDATA_int[25]));

	qlIBUF QL_INST_A2F_L_11_2 (.IN_IBUF(lint_WDATA[26]),.OUT_IBUF(lint_WDATA_int[26]));

	qlIBUF QL_INST_A2F_L_11_3 (.IN_IBUF(lint_WDATA[27]),.OUT_IBUF(lint_WDATA_int[27]));

	qlIBUF QL_INST_A2F_L_11_4 (.IN_IBUF(lint_WDATA[28]),.OUT_IBUF(lint_WDATA_int[28]));

	qlIBUF QL_INST_A2F_L_11_5 (.IN_IBUF(lint_WDATA[29]),.OUT_IBUF(lint_WDATA_int[29]));

	qlOBUF QL_INST_F2A_L_12_8 (.IN_OBUF(lint_RDATA_dup_0[0]),.OUT_OBUF(lint_RDATA[0]));

	qlOBUF QL_INST_F2A_L_12_9 (.IN_OBUF(lint_RDATA_dup_0[1]),.OUT_OBUF(lint_RDATA[1]));

	qlOBUF QL_INST_F2A_L_12_10 (.IN_OBUF(lint_RDATA_dup_0[2]),.OUT_OBUF(lint_RDATA[2]));

	qlOBUF QL_INST_F2A_L_12_11 (.IN_OBUF(lint_RDATA_dup_0[3]),.OUT_OBUF(lint_RDATA[3]));

	qlOBUF QL_INST_F2A_L_12_12 (.IN_OBUF(lint_RDATA_dup_0[4]),.OUT_OBUF(lint_RDATA[4]));

	qlOBUF QL_INST_F2A_L_12_13 (.IN_OBUF(lint_RDATA_dup_0[5]),.OUT_OBUF(lint_RDATA[5]));

	qlOBUF QL_INST_F2A_L_12_14 (.IN_OBUF(lint_RDATA_dup_0[6]),.OUT_OBUF(lint_RDATA[6]));

	qlOBUF QL_INST_F2A_L_12_15 (.IN_OBUF(lint_RDATA_dup_0[7]),.OUT_OBUF(lint_RDATA[7]));

	qlOBUF QL_INST_F2A_L_12_16 (.IN_OBUF(lint_RDATA_dup_0[8]),.OUT_OBUF(lint_RDATA[8]));

	qlIBUF QL_INST_A2F_L_12_0 (.IN_IBUF(lint_WDATA[30]),.OUT_IBUF(lint_WDATA_int[30]));

	qlIBUF QL_INST_A2F_L_12_1 (.IN_IBUF(lint_WDATA[31]),.OUT_IBUF(lint_WDATA_int[31]));

	qlIBUF QL_INST_A2F_L_12_2 (.IN_IBUF(lint_REQ),.OUT_IBUF(lint_REQ_int));

	qlIBUF QL_INST_A2F_L_12_3 (.IN_IBUF(lint_WEN),.OUT_IBUF(lint_WEN_int));

	qlIBUF QL_INST_A2F_L_12_4 (.IN_IBUF(lint_BE[0]),.OUT_IBUF(lint_BE_int[0]));

	qlIBUF QL_INST_A2F_L_12_5 (.IN_IBUF(lint_BE[1]),.OUT_IBUF(lint_BE_int[1]));

	qlIBUF QL_INST_A2F_L_12_6 (.IN_IBUF(lint_BE[2]),.OUT_IBUF(lint_BE_int[2]));

	qlIBUF QL_INST_A2F_L_12_7 (.IN_IBUF(lint_BE[3]),.OUT_IBUF(lint_BE_int[3]));

	qlOBUF QL_INST_F2A_L_13_0 (.IN_OBUF(lint_RDATA_dup_0[9]),.OUT_OBUF(lint_RDATA[9]));

	qlOBUF QL_INST_F2A_L_13_1 (.IN_OBUF(lint_RDATA_dup_0[10]),.OUT_OBUF(lint_RDATA[10]));

	qlOBUF QL_INST_F2A_L_13_2 (.IN_OBUF(lint_RDATA_dup_0[11]),.OUT_OBUF(lint_RDATA[11]));

	qlOBUF QL_INST_F2A_L_13_3 (.IN_OBUF(lint_RDATA_dup_0[12]),.OUT_OBUF(lint_RDATA[12]));

	qlOBUF QL_INST_F2A_L_13_4 (.IN_OBUF(lint_RDATA_dup_0[13]),.OUT_OBUF(lint_RDATA[13]));

	qlOBUF QL_INST_F2A_L_13_5 (.IN_OBUF(lint_RDATA_dup_0[14]),.OUT_OBUF(lint_RDATA[14]));

	qlOBUF QL_INST_F2A_L_13_6 (.IN_OBUF(lint_RDATA_dup_0[15]),.OUT_OBUF(lint_RDATA[15]));

	qlIBUF QL_INST_A2F_L_13_0 (.IN_IBUF(lint_ADDR[0]),.OUT_IBUF(lint_ADDR_int[0]));

	qlIBUF QL_INST_A2F_L_13_1 (.IN_IBUF(lint_ADDR[1]),.OUT_IBUF(lint_ADDR_int[1]));

	qlIBUF QL_INST_A2F_L_13_2 (.IN_IBUF(lint_ADDR[2]),.OUT_IBUF(lint_ADDR_int[2]));

	qlIBUF QL_INST_A2F_L_13_3 (.IN_IBUF(lint_ADDR[3]),.OUT_IBUF(lint_ADDR_int[3]));

	qlIBUF QL_INST_A2F_L_13_4 (.IN_IBUF(lint_ADDR[4]),.OUT_IBUF(lint_ADDR_int[4]));

	qlIBUF QL_INST_A2F_L_13_5 (.IN_IBUF(lint_ADDR[5]),.OUT_IBUF(lint_ADDR_int[5]));

	qlOBUF QL_INST_F2A_L_14_0 (.IN_OBUF(CLK_int_0__CAND0_TLSBL_0_padClk),.OUT_OBUF(lint_clk));

	qlOBUF QL_INST_F2A_L_14_1 (.IN_OBUF(lint_RDATA_dup_0[16]),.OUT_OBUF(lint_RDATA[16]));

	qlOBUF QL_INST_F2A_L_14_2 (.IN_OBUF(lint_RDATA_dup_0[17]),.OUT_OBUF(lint_RDATA[17]));

	qlOBUF QL_INST_F2A_L_14_3 (.IN_OBUF(lint_RDATA_dup_0[18]),.OUT_OBUF(lint_RDATA[18]));

	qlOBUF QL_INST_F2A_L_14_4 (.IN_OBUF(lint_RDATA_dup_0[19]),.OUT_OBUF(lint_RDATA[19]));

	qlOBUF QL_INST_F2A_L_14_5 (.IN_OBUF(lint_RDATA_dup_0[20]),.OUT_OBUF(lint_RDATA[20]));

	qlOBUF QL_INST_F2A_L_14_6 (.IN_OBUF(lint_RDATA_dup_0[21]),.OUT_OBUF(lint_RDATA[21]));

	qlOBUF QL_INST_F2A_L_14_7 (.IN_OBUF(lint_RDATA_dup_0[22]),.OUT_OBUF(lint_RDATA[22]));

	qlOBUF QL_INST_F2A_L_14_8 (.IN_OBUF(lint_RDATA_dup_0[23]),.OUT_OBUF(lint_RDATA[23]));

	qlOBUF QL_INST_F2A_L_14_9 (.IN_OBUF(lint_VALID_dup_0),.OUT_OBUF(lint_VALID));

	qlIBUF QL_INST_A2F_L_14_0 (.IN_IBUF(lint_ADDR[6]),.OUT_IBUF(lint_ADDR_int[6]));

	qlIBUF QL_INST_A2F_L_14_1 (.IN_IBUF(lint_ADDR[7]),.OUT_IBUF(lint_ADDR_int[7]));

	qlIBUF QL_INST_A2F_L_14_2 (.IN_IBUF(lint_ADDR[8]),.OUT_IBUF(lint_ADDR_int[8]));

	qlIBUF QL_INST_A2F_L_14_3 (.IN_IBUF(lint_ADDR[9]),.OUT_IBUF(lint_ADDR_int[9]));

	qlIBUF QL_INST_A2F_L_14_4 (.IN_IBUF(lint_ADDR[10]),.OUT_IBUF(lint_ADDR_int[10]));

	qlIBUF QL_INST_A2F_L_14_5 (.IN_IBUF(lint_ADDR[11]),.OUT_IBUF(lint_ADDR_int[11]));

	qlIBUF QL_INST_A2F_L_14_6 (.IN_IBUF(lint_ADDR[12]),.OUT_IBUF(lint_ADDR_int[12]));

	qlIBUF QL_INST_A2F_L_14_7 (.IN_IBUF(lint_ADDR[13]),.OUT_IBUF(lint_ADDR_int[13]));

	qlOBUF QL_INST_F2A_L_15_0 (.IN_OBUF(lint_RDATA_dup_0[24]),.OUT_OBUF(lint_RDATA[24]));

	qlOBUF QL_INST_F2A_L_15_1 (.IN_OBUF(lint_RDATA_dup_0[25]),.OUT_OBUF(lint_RDATA[25]));

	qlOBUF QL_INST_F2A_L_15_2 (.IN_OBUF(lint_RDATA_dup_0[26]),.OUT_OBUF(lint_RDATA[26]));

	qlOBUF QL_INST_F2A_L_15_3 (.IN_OBUF(lint_RDATA_dup_0[27]),.OUT_OBUF(lint_RDATA[27]));

	qlOBUF QL_INST_F2A_L_15_4 (.IN_OBUF(lint_RDATA_dup_0[28]),.OUT_OBUF(lint_RDATA[28]));

	qlOBUF QL_INST_F2A_L_15_5 (.IN_OBUF(lint_RDATA_dup_0[29]),.OUT_OBUF(lint_RDATA[29]));

	qlOBUF QL_INST_F2A_L_15_6 (.IN_OBUF(lint_RDATA_dup_0[30]),.OUT_OBUF(lint_RDATA[30]));

	qlOBUF QL_INST_F2A_L_15_7 (.IN_OBUF(lint_RDATA_dup_0[31]),.OUT_OBUF(lint_RDATA[31]));

	qlOBUF QL_INST_F2A_L_15_8 (.IN_OBUF(lint_GNT_dup_0),.OUT_OBUF(lint_GNT));

	qlIBUF QL_INST_A2F_L_15_0 (.IN_IBUF(lint_ADDR[14]),.OUT_IBUF(lint_ADDR_int[14]));

	qlIBUF QL_INST_A2F_L_15_1 (.IN_IBUF(lint_ADDR[15]),.OUT_IBUF(lint_ADDR_int[15]));

	qlIBUF QL_INST_A2F_L_15_2 (.IN_IBUF(lint_ADDR[16]),.OUT_IBUF(lint_ADDR_int[16]));

	qlIBUF QL_INST_A2F_L_15_3 (.IN_IBUF(lint_ADDR[17]),.OUT_IBUF(lint_ADDR_int[17]));

	qlIBUF QL_INST_A2F_L_15_4 (.IN_IBUF(lint_ADDR[18]),.OUT_IBUF(lint_ADDR_int[18]));

	qlIBUF QL_INST_A2F_L_15_5 (.IN_IBUF(lint_ADDR[19]),.OUT_IBUF(lint_ADDR_int[19]));

	qlIBUF QL_INST_A2F_L_16_0 (.IN_IBUF(fpgaio_in[64]),.OUT_IBUF(fpgaio_in_int[64]));

	qlIBUF QL_INST_A2F_L_16_1 (.IN_IBUF(fpgaio_in[65]),.OUT_IBUF(fpgaio_in_int[65]));

	qlIBUF QL_INST_A2F_L_16_2 (.IN_IBUF(fpgaio_in[66]),.OUT_IBUF(fpgaio_in_int[66]));

	qlIBUF QL_INST_A2F_L_16_3 (.IN_IBUF(fpgaio_in[67]),.OUT_IBUF(fpgaio_in_int[67]));

	qlIBUF QL_INST_A2F_L_16_4 (.IN_IBUF(fpgaio_in[68]),.OUT_IBUF(fpgaio_in_int[68]));

	qlIBUF QL_INST_A2F_L_16_5 (.IN_IBUF(fpgaio_in[69]),.OUT_IBUF(fpgaio_in_int[69]));

	qlIBUF QL_INST_A2F_L_16_6 (.IN_IBUF(fpgaio_in[70]),.OUT_IBUF(fpgaio_in_int[70]));

	qlIBUF QL_INST_A2F_L_16_7 (.IN_IBUF(fpgaio_in[71]),.OUT_IBUF(fpgaio_in_int[71]));

	qlOBUF QL_INST_F2A_L_17_0 (.IN_OBUF(fpgaio_out_dup_0[64]),.OUT_OBUF(fpgaio_out[64]));

	qlOBUF QL_INST_F2A_L_17_1 (.IN_OBUF(fpgaio_oe_dup_0[64]),.OUT_OBUF(fpgaio_oe[64]));

	qlOBUF QL_INST_F2A_L_17_2 (.IN_OBUF(fpgaio_out_dup_0[65]),.OUT_OBUF(fpgaio_out[65]));

	qlOBUF QL_INST_F2A_L_17_3 (.IN_OBUF(fpgaio_oe_dup_0[65]),.OUT_OBUF(fpgaio_oe[65]));

	qlOBUF QL_INST_F2A_L_17_4 (.IN_OBUF(fpgaio_out_dup_0[66]),.OUT_OBUF(fpgaio_out[66]));

	qlOBUF QL_INST_F2A_L_17_5 (.IN_OBUF(fpgaio_oe_dup_0[66]),.OUT_OBUF(fpgaio_oe[66]));

	qlOBUF QL_INST_F2A_L_17_6 (.IN_OBUF(fpgaio_out_dup_0[67]),.OUT_OBUF(fpgaio_out[67]));

	qlOBUF QL_INST_F2A_L_17_7 (.IN_OBUF(fpgaio_oe_dup_0[67]),.OUT_OBUF(fpgaio_oe[67]));

	qlIBUF QL_INST_A2F_L_17_0 (.IN_IBUF(fpgaio_in[72]),.OUT_IBUF(fpgaio_in_int[72]));

	qlIBUF QL_INST_A2F_L_17_1 (.IN_IBUF(fpgaio_in[73]),.OUT_IBUF(fpgaio_in_int[73]));

	qlIBUF QL_INST_A2F_L_17_2 (.IN_IBUF(fpgaio_in[74]),.OUT_IBUF(fpgaio_in_int[74]));

	qlIBUF QL_INST_A2F_L_17_3 (.IN_IBUF(fpgaio_in[75]),.OUT_IBUF(fpgaio_in_int[75]));

	qlIBUF QL_INST_A2F_L_17_4 (.IN_IBUF(fpgaio_in[76]),.OUT_IBUF(fpgaio_in_int[76]));

	qlIBUF QL_INST_A2F_L_17_5 (.IN_IBUF(fpgaio_in[77]),.OUT_IBUF(fpgaio_in_int[77]));

	qlOBUF QL_INST_F2A_L_18_0 (.IN_OBUF(fpgaio_out_dup_0[68]),.OUT_OBUF(fpgaio_out[68]));

	qlOBUF QL_INST_F2A_L_18_1 (.IN_OBUF(fpgaio_oe_dup_0[68]),.OUT_OBUF(fpgaio_oe[68]));

	qlOBUF QL_INST_F2A_L_18_2 (.IN_OBUF(fpgaio_out_dup_0[69]),.OUT_OBUF(fpgaio_out[69]));

	qlOBUF QL_INST_F2A_L_18_3 (.IN_OBUF(fpgaio_oe_dup_0[69]),.OUT_OBUF(fpgaio_oe[69]));

	qlOBUF QL_INST_F2A_L_18_4 (.IN_OBUF(fpgaio_out_dup_0[70]),.OUT_OBUF(fpgaio_out[70]));

	qlOBUF QL_INST_F2A_L_18_5 (.IN_OBUF(fpgaio_oe_dup_0[70]),.OUT_OBUF(fpgaio_oe[70]));

	qlOBUF QL_INST_F2A_L_18_6 (.IN_OBUF(fpgaio_out_dup_0[71]),.OUT_OBUF(fpgaio_out[71]));

	qlOBUF QL_INST_F2A_L_18_7 (.IN_OBUF(fpgaio_oe_dup_0[71]),.OUT_OBUF(fpgaio_oe[71]));

	qlOBUF QL_INST_F2A_L_18_8 (.IN_OBUF(fpgaio_out_dup_0[72]),.OUT_OBUF(fpgaio_out[72]));

	qlOBUF QL_INST_F2A_L_18_9 (.IN_OBUF(fpgaio_oe_dup_0[72]),.OUT_OBUF(fpgaio_oe[72]));

	qlOBUF QL_INST_F2A_L_18_10 (.IN_OBUF(fpgaio_out_dup_0[73]),.OUT_OBUF(fpgaio_out[73]));

	qlOBUF QL_INST_F2A_L_18_11 (.IN_OBUF(fpgaio_oe_dup_0[73]),.OUT_OBUF(fpgaio_oe[73]));

	qlOBUF QL_INST_F2A_L_18_12 (.IN_OBUF(fpgaio_out_dup_0[74]),.OUT_OBUF(fpgaio_out[74]));

	qlOBUF QL_INST_F2A_L_18_13 (.IN_OBUF(fpgaio_oe_dup_0[74]),.OUT_OBUF(fpgaio_oe[74]));

	qlOBUF QL_INST_F2A_L_18_14 (.IN_OBUF(fpgaio_out_dup_0[75]),.OUT_OBUF(fpgaio_out[75]));

	qlOBUF QL_INST_F2A_L_18_15 (.IN_OBUF(fpgaio_oe_dup_0[75]),.OUT_OBUF(fpgaio_oe[75]));

	qlIBUF QL_INST_A2F_L_18_0 (.IN_IBUF(fpgaio_in[78]),.OUT_IBUF(fpgaio_in_int[78]));

	qlIBUF QL_INST_A2F_L_18_1 (.IN_IBUF(fpgaio_in[79]),.OUT_IBUF(fpgaio_in_int[79]));

	qlOBUF QL_INST_F2A_L_19_0 (.IN_OBUF(fpgaio_out_dup_0[76]),.OUT_OBUF(fpgaio_out[76]));

	qlOBUF QL_INST_F2A_L_19_1 (.IN_OBUF(fpgaio_oe_dup_0[76]),.OUT_OBUF(fpgaio_oe[76]));

	qlOBUF QL_INST_F2A_L_19_2 (.IN_OBUF(fpgaio_out_dup_0[77]),.OUT_OBUF(fpgaio_out[77]));

	qlOBUF QL_INST_F2A_L_19_3 (.IN_OBUF(fpgaio_oe_dup_0[77]),.OUT_OBUF(fpgaio_oe[77]));

	qlOBUF QL_INST_F2A_L_19_4 (.IN_OBUF(fpgaio_out_dup_0[78]),.OUT_OBUF(fpgaio_out[78]));

	qlOBUF QL_INST_F2A_L_19_5 (.IN_OBUF(fpgaio_oe_dup_0[78]),.OUT_OBUF(fpgaio_oe[78]));

	qlOBUF QL_INST_F2A_L_19_6 (.IN_OBUF(fpgaio_out_dup_0[79]),.OUT_OBUF(fpgaio_out[79]));

	qlOBUF QL_INST_F2A_L_19_7 (.IN_OBUF(fpgaio_oe_dup_0[79]),.OUT_OBUF(fpgaio_oe[79]));

	qlIBUF QL_INST_A2F_L_19_0 (.IN_IBUF(control_in[0]),.OUT_IBUF(control_in_int[0]));

	qlIBUF QL_INST_A2F_L_19_1 (.IN_IBUF(control_in[1]),.OUT_IBUF(control_in_int[1]));

	qlIBUF QL_INST_A2F_L_19_2 (.IN_IBUF(control_in[2]),.OUT_IBUF(control_in_int[2]));

	qlIBUF QL_INST_A2F_L_19_3 (.IN_IBUF(control_in[3]),.OUT_IBUF(control_in_int[3]));

	qlIBUF QL_INST_A2F_L_19_4 (.IN_IBUF(control_in[4]),.OUT_IBUF(control_in_int[4]));

	qlIBUF QL_INST_A2F_L_19_5 (.IN_IBUF(control_in[5]),.OUT_IBUF(control_in_int[5]));

	qlOBUF QL_INST_F2A_L_20_0 (.IN_OBUF(control_in_int[0]),.OUT_OBUF(status_out[0]));

	qlOBUF QL_INST_F2A_L_20_1 (.IN_OBUF(control_in_int[1]),.OUT_OBUF(status_out[1]));

	qlOBUF QL_INST_F2A_L_20_2 (.IN_OBUF(control_in_int[2]),.OUT_OBUF(status_out[2]));

	qlOBUF QL_INST_F2A_L_20_3 (.IN_OBUF(control_in_int[3]),.OUT_OBUF(status_out[3]));

	qlOBUF QL_INST_F2A_L_20_4 (.IN_OBUF(control_in_int[4]),.OUT_OBUF(status_out[4]));

	qlOBUF QL_INST_F2A_L_20_5 (.IN_OBUF(control_in_int[5]),.OUT_OBUF(status_out[5]));

	qlOBUF QL_INST_F2A_L_20_6 (.IN_OBUF(control_in_int[6]),.OUT_OBUF(status_out[6]));

	qlOBUF QL_INST_F2A_L_20_7 (.IN_OBUF(control_in_int[7]),.OUT_OBUF(status_out[7]));

	qlOBUF QL_INST_F2A_L_20_8 (.IN_OBUF(control_in_int[8]),.OUT_OBUF(status_out[8]));

	qlOBUF QL_INST_F2A_L_20_9 (.IN_OBUF(control_in_int[9]),.OUT_OBUF(status_out[9]));

	qlOBUF QL_INST_F2A_L_20_10 (.IN_OBUF(control_in_int[10]),.OUT_OBUF(status_out[10]));

	qlOBUF QL_INST_F2A_L_20_11 (.IN_OBUF(control_in_int[11]),.OUT_OBUF(status_out[11]));

	qlOBUF QL_INST_F2A_L_20_12 (.IN_OBUF(control_in_int[12]),.OUT_OBUF(status_out[12]));

	qlOBUF QL_INST_F2A_L_20_13 (.IN_OBUF(control_in_int[13]),.OUT_OBUF(status_out[13]));

	qlOBUF QL_INST_F2A_L_20_14 (.IN_OBUF(control_in_int[14]),.OUT_OBUF(status_out[14]));

	qlOBUF QL_INST_F2A_L_20_15 (.IN_OBUF(control_in_int[15]),.OUT_OBUF(status_out[15]));

	qlOBUF QL_INST_F2A_L_20_16 (.IN_OBUF(control_in_int[16]),.OUT_OBUF(status_out[16]));

	qlOBUF QL_INST_F2A_L_20_17 (.IN_OBUF(control_in_int[17]),.OUT_OBUF(status_out[17]));

	qlIBUF QL_INST_A2F_L_20_0 (.IN_IBUF(control_in[6]),.OUT_IBUF(control_in_int[6]));

	qlIBUF QL_INST_A2F_L_20_1 (.IN_IBUF(control_in[7]),.OUT_IBUF(control_in_int[7]));

	qlIBUF QL_INST_A2F_L_20_2 (.IN_IBUF(control_in[8]),.OUT_IBUF(control_in_int[8]));

	qlIBUF QL_INST_A2F_L_20_3 (.IN_IBUF(control_in[9]),.OUT_IBUF(control_in_int[9]));

	qlIBUF QL_INST_A2F_L_20_4 (.IN_IBUF(control_in[10]),.OUT_IBUF(control_in_int[10]));

	qlIBUF QL_INST_A2F_L_20_5 (.IN_IBUF(control_in[11]),.OUT_IBUF(control_in_int[11]));

	qlIBUF QL_INST_A2F_L_20_6 (.IN_IBUF(control_in[12]),.OUT_IBUF(control_in_int[12]));

	qlIBUF QL_INST_A2F_L_20_7 (.IN_IBUF(control_in[13]),.OUT_IBUF(control_in_int[13]));

	qlOBUF QL_INST_F2A_L_21_0 (.IN_OBUF(control_in_int[18]),.OUT_OBUF(status_out[18]));

	qlOBUF QL_INST_F2A_L_21_1 (.IN_OBUF(control_in_int[19]),.OUT_OBUF(status_out[19]));

	qlOBUF QL_INST_F2A_L_21_2 (.IN_OBUF(control_in_int[20]),.OUT_OBUF(status_out[20]));

	qlOBUF QL_INST_F2A_L_21_3 (.IN_OBUF(control_in_int[21]),.OUT_OBUF(status_out[21]));

	qlOBUF QL_INST_F2A_L_21_4 (.IN_OBUF(control_in_int[22]),.OUT_OBUF(status_out[22]));

	qlOBUF QL_INST_F2A_L_21_5 (.IN_OBUF(control_in_int[23]),.OUT_OBUF(status_out[23]));

	qlOBUF QL_INST_F2A_L_21_6 (.IN_OBUF(control_in_int[24]),.OUT_OBUF(status_out[24]));

	qlOBUF QL_INST_F2A_L_21_7 (.IN_OBUF(control_in_int[25]),.OUT_OBUF(status_out[25]));

	qlOBUF QL_INST_F2A_L_21_8 (.IN_OBUF(control_in_int[26]),.OUT_OBUF(status_out[26]));

	qlOBUF QL_INST_F2A_L_21_9 (.IN_OBUF(control_in_int[27]),.OUT_OBUF(status_out[27]));

	qlOBUF QL_INST_F2A_L_21_10 (.IN_OBUF(control_in_int[28]),.OUT_OBUF(status_out[28]));

	qlOBUF QL_INST_F2A_L_21_11 (.IN_OBUF(control_in_int[29]),.OUT_OBUF(status_out[29]));

	qlIBUF QL_INST_A2F_L_21_0 (.IN_IBUF(control_in[14]),.OUT_IBUF(control_in_int[14]));

	qlIBUF QL_INST_A2F_L_21_1 (.IN_IBUF(control_in[15]),.OUT_IBUF(control_in_int[15]));

	qlIBUF QL_INST_A2F_L_21_2 (.IN_IBUF(control_in[16]),.OUT_IBUF(control_in_int[16]));

	qlIBUF QL_INST_A2F_L_21_3 (.IN_IBUF(control_in[17]),.OUT_IBUF(control_in_int[17]));

	qlIBUF QL_INST_A2F_L_21_4 (.IN_IBUF(control_in[18]),.OUT_IBUF(control_in_int[18]));

	qlIBUF QL_INST_A2F_L_21_5 (.IN_IBUF(control_in[19]),.OUT_IBUF(control_in_int[19]));

	qlOBUF QL_INST_F2A_L_22_0 (.IN_OBUF(control_in_int[30]),.OUT_OBUF(status_out[30]));

	qlOBUF QL_INST_F2A_L_22_1 (.IN_OBUF(control_in_int[31]),.OUT_OBUF(status_out[31]));

	qlIBUF QL_INST_A2F_L_22_0 (.IN_IBUF(control_in[20]),.OUT_IBUF(control_in_int[20]));

	qlIBUF QL_INST_A2F_L_22_1 (.IN_IBUF(control_in[21]),.OUT_IBUF(control_in_int[21]));

	qlIBUF QL_INST_A2F_L_22_2 (.IN_IBUF(control_in[22]),.OUT_IBUF(control_in_int[22]));

	qlIBUF QL_INST_A2F_L_22_3 (.IN_IBUF(control_in[23]),.OUT_IBUF(control_in_int[23]));

	qlIBUF QL_INST_A2F_L_22_4 (.IN_IBUF(control_in[24]),.OUT_IBUF(control_in_int[24]));

	qlIBUF QL_INST_A2F_L_22_5 (.IN_IBUF(control_in[25]),.OUT_IBUF(control_in_int[25]));

	qlIBUF QL_INST_A2F_L_22_6 (.IN_IBUF(control_in[26]),.OUT_IBUF(control_in_int[26]));

	qlIBUF QL_INST_A2F_L_23_0 (.IN_IBUF(control_in[27]),.OUT_IBUF(control_in_int[27]));

	qlIBUF QL_INST_A2F_L_23_1 (.IN_IBUF(control_in[28]),.OUT_IBUF(control_in_int[28]));

	qlIBUF QL_INST_A2F_L_23_2 (.IN_IBUF(control_in[29]),.OUT_IBUF(control_in_int[29]));

	qlIBUF QL_INST_A2F_L_23_3 (.IN_IBUF(control_in[30]),.OUT_IBUF(control_in_int[30]));

	qlIBUF QL_INST_A2F_L_23_4 (.IN_IBUF(control_in[31]),.OUT_IBUF(control_in_int[31]));

	qlOBUF QL_INST_F2A_L_25_0 (.IN_OBUF(fpgaio_out_dup_0[32]),.OUT_OBUF(fpgaio_out[32]));

	qlOBUF QL_INST_F2A_L_25_1 (.IN_OBUF(fpgaio_oe_dup_0[32]),.OUT_OBUF(fpgaio_oe[32]));

	qlOBUF QL_INST_F2A_L_25_2 (.IN_OBUF(fpgaio_out_dup_0[33]),.OUT_OBUF(fpgaio_out[33]));

	qlOBUF QL_INST_F2A_L_25_3 (.IN_OBUF(fpgaio_oe_dup_0[33]),.OUT_OBUF(fpgaio_oe[33]));

	qlOBUF QL_INST_F2A_L_25_4 (.IN_OBUF(fpgaio_out_dup_0[34]),.OUT_OBUF(fpgaio_out[34]));

	qlOBUF QL_INST_F2A_L_25_5 (.IN_OBUF(fpgaio_oe_dup_0[34]),.OUT_OBUF(fpgaio_oe[34]));

	qlOBUF QL_INST_F2A_L_25_6 (.IN_OBUF(fpgaio_out_dup_0[35]),.OUT_OBUF(fpgaio_out[35]));

	qlOBUF QL_INST_F2A_L_25_7 (.IN_OBUF(fpgaio_oe_dup_0[35]),.OUT_OBUF(fpgaio_oe[35]));

	qlOBUF QL_INST_F2A_L_25_8 (.IN_OBUF(fpgaio_in_int[8]),.OUT_OBUF(events_o[8]));

	qlIBUF QL_INST_A2F_L_25_0 (.IN_IBUF(fpgaio_in[32]),.OUT_IBUF(fpgaio_in_int[32]));

	qlIBUF QL_INST_A2F_L_25_1 (.IN_IBUF(fpgaio_in[33]),.OUT_IBUF(fpgaio_in_int[33]));

	qlIBUF QL_INST_A2F_L_25_2 (.IN_IBUF(RESET[2]),.OUT_IBUF(RESET_int[2]));

	qlIBUF QL_INST_A2F_L_25_3 (.IN_IBUF(fpgaio_in[34]),.OUT_IBUF(fpgaio_in_int[34]));

	qlIBUF QL_INST_A2F_L_25_4 (.IN_IBUF(fpgaio_in[35]),.OUT_IBUF(fpgaio_in_int[35]));

	qlOBUF QL_INST_F2A_L_26_0 (.IN_OBUF(fpgaio_out_dup_0[36]),.OUT_OBUF(fpgaio_out[36]));

	qlOBUF QL_INST_F2A_L_26_1 (.IN_OBUF(fpgaio_oe_dup_0[36]),.OUT_OBUF(fpgaio_oe[36]));

	qlOBUF QL_INST_F2A_L_26_2 (.IN_OBUF(fpgaio_out_dup_0[37]),.OUT_OBUF(fpgaio_out[37]));

	qlOBUF QL_INST_F2A_L_26_3 (.IN_OBUF(fpgaio_oe_dup_0[37]),.OUT_OBUF(fpgaio_oe[37]));

	qlOBUF QL_INST_F2A_L_26_4 (.IN_OBUF(fpgaio_out_dup_0[38]),.OUT_OBUF(fpgaio_out[38]));

	qlOBUF QL_INST_F2A_L_26_5 (.IN_OBUF(fpgaio_oe_dup_0[38]),.OUT_OBUF(fpgaio_oe[38]));

	qlOBUF QL_INST_F2A_L_26_6 (.IN_OBUF(fpgaio_out_dup_0[39]),.OUT_OBUF(fpgaio_out[39]));

	qlOBUF QL_INST_F2A_L_26_7 (.IN_OBUF(fpgaio_oe_dup_0[39]),.OUT_OBUF(fpgaio_oe[39]));

	qlOBUF QL_INST_F2A_L_26_8 (.IN_OBUF(fpgaio_in_int[9]),.OUT_OBUF(events_o[9]));

	qlIBUF QL_INST_A2F_L_26_0 (.IN_IBUF(fpgaio_in[36]),.OUT_IBUF(fpgaio_in_int[36]));

	qlIBUF QL_INST_A2F_L_26_1 (.IN_IBUF(fpgaio_in[37]),.OUT_IBUF(fpgaio_in_int[37]));

	qlIBUF QL_INST_A2F_L_26_2 (.IN_IBUF(fpgaio_in[38]),.OUT_IBUF(fpgaio_in_int[38]));

	qlIBUF QL_INST_A2F_L_26_3 (.IN_IBUF(fpgaio_in[39]),.OUT_IBUF(fpgaio_in_int[39]));

	qlOBUF QL_INST_F2A_L_27_0 (.IN_OBUF(fpgaio_out_dup_0[40]),.OUT_OBUF(fpgaio_out[40]));

	qlOBUF QL_INST_F2A_L_27_1 (.IN_OBUF(fpgaio_oe_dup_0[40]),.OUT_OBUF(fpgaio_oe[40]));

	qlOBUF QL_INST_F2A_L_27_2 (.IN_OBUF(fpgaio_out_dup_0[41]),.OUT_OBUF(fpgaio_out[41]));

	qlOBUF QL_INST_F2A_L_27_3 (.IN_OBUF(fpgaio_oe_dup_0[41]),.OUT_OBUF(fpgaio_oe[41]));

	qlOBUF QL_INST_F2A_L_27_4 (.IN_OBUF(fpgaio_out_dup_0[42]),.OUT_OBUF(fpgaio_out[42]));

	qlOBUF QL_INST_F2A_L_27_5 (.IN_OBUF(fpgaio_oe_dup_0[42]),.OUT_OBUF(fpgaio_oe[42]));

	qlOBUF QL_INST_F2A_L_27_6 (.IN_OBUF(fpgaio_out_dup_0[43]),.OUT_OBUF(fpgaio_out[43]));

	qlOBUF QL_INST_F2A_L_27_7 (.IN_OBUF(fpgaio_oe_dup_0[43]),.OUT_OBUF(fpgaio_oe[43]));

	qlOBUF QL_INST_F2A_L_27_8 (.IN_OBUF(fpgaio_in_int[10]),.OUT_OBUF(events_o[10]));

	qlIBUF QL_INST_A2F_L_27_0 (.IN_IBUF(fpgaio_in[40]),.OUT_IBUF(fpgaio_in_int[40]));

	qlIBUF QL_INST_A2F_L_27_1 (.IN_IBUF(fpgaio_in[41]),.OUT_IBUF(fpgaio_in_int[41]));

	qlIBUF QL_INST_A2F_L_27_2 (.IN_IBUF(fpgaio_in[42]),.OUT_IBUF(fpgaio_in_int[42]));

	qlIBUF QL_INST_A2F_L_27_3 (.IN_IBUF(fpgaio_in[43]),.OUT_IBUF(fpgaio_in_int[43]));

	qlOBUF QL_INST_F2A_L_28_0 (.IN_OBUF(fpgaio_out_dup_0[44]),.OUT_OBUF(fpgaio_out[44]));

	qlOBUF QL_INST_F2A_L_28_1 (.IN_OBUF(fpgaio_oe_dup_0[44]),.OUT_OBUF(fpgaio_oe[44]));

	qlOBUF QL_INST_F2A_L_28_2 (.IN_OBUF(fpgaio_out_dup_0[45]),.OUT_OBUF(fpgaio_out[45]));

	qlOBUF QL_INST_F2A_L_28_3 (.IN_OBUF(fpgaio_oe_dup_0[45]),.OUT_OBUF(fpgaio_oe[45]));

	qlOBUF QL_INST_F2A_L_28_4 (.IN_OBUF(fpgaio_out_dup_0[46]),.OUT_OBUF(fpgaio_out[46]));

	qlOBUF QL_INST_F2A_L_28_5 (.IN_OBUF(fpgaio_oe_dup_0[46]),.OUT_OBUF(fpgaio_oe[46]));

	qlOBUF QL_INST_F2A_L_28_6 (.IN_OBUF(fpgaio_out_dup_0[47]),.OUT_OBUF(fpgaio_out[47]));

	qlOBUF QL_INST_F2A_L_28_7 (.IN_OBUF(fpgaio_oe_dup_0[47]),.OUT_OBUF(fpgaio_oe[47]));

	qlOBUF QL_INST_F2A_L_28_8 (.IN_OBUF(fpgaio_in_int[11]),.OUT_OBUF(events_o[11]));

	qlIBUF QL_INST_A2F_L_28_0 (.IN_IBUF(fpgaio_in[44]),.OUT_IBUF(fpgaio_in_int[44]));

	qlIBUF QL_INST_A2F_L_28_1 (.IN_IBUF(fpgaio_in[45]),.OUT_IBUF(fpgaio_in_int[45]));

	qlIBUF QL_INST_A2F_L_28_2 (.IN_IBUF(fpgaio_in[46]),.OUT_IBUF(fpgaio_in_int[46]));

	qlIBUF QL_INST_A2F_L_28_3 (.IN_IBUF(fpgaio_in[47]),.OUT_IBUF(fpgaio_in_int[47]));

	qlOBUF QL_INST_F2A_L_29_0 (.IN_OBUF(fpgaio_out_dup_0[48]),.OUT_OBUF(fpgaio_out[48]));

	qlOBUF QL_INST_F2A_L_29_1 (.IN_OBUF(fpgaio_oe_dup_0[48]),.OUT_OBUF(fpgaio_oe[48]));

	qlOBUF QL_INST_F2A_L_29_2 (.IN_OBUF(fpgaio_out_dup_0[49]),.OUT_OBUF(fpgaio_out[49]));

	qlOBUF QL_INST_F2A_L_29_3 (.IN_OBUF(fpgaio_oe_dup_0[49]),.OUT_OBUF(fpgaio_oe[49]));

	qlOBUF QL_INST_F2A_L_29_4 (.IN_OBUF(fpgaio_out_dup_0[50]),.OUT_OBUF(fpgaio_out[50]));

	qlOBUF QL_INST_F2A_L_29_5 (.IN_OBUF(fpgaio_oe_dup_0[50]),.OUT_OBUF(fpgaio_oe[50]));

	qlOBUF QL_INST_F2A_L_29_6 (.IN_OBUF(fpgaio_out_dup_0[51]),.OUT_OBUF(fpgaio_out[51]));

	qlOBUF QL_INST_F2A_L_29_7 (.IN_OBUF(fpgaio_oe_dup_0[51]),.OUT_OBUF(fpgaio_oe[51]));

	qlOBUF QL_INST_F2A_L_29_8 (.IN_OBUF(fpgaio_in_int[12]),.OUT_OBUF(events_o[12]));

	qlIBUF QL_INST_A2F_L_29_0 (.IN_IBUF(fpgaio_in[48]),.OUT_IBUF(fpgaio_in_int[48]));

	qlIBUF QL_INST_A2F_L_29_1 (.IN_IBUF(fpgaio_in[49]),.OUT_IBUF(fpgaio_in_int[49]));

	qlIBUF QL_INST_A2F_L_29_2 (.IN_IBUF(fpgaio_in[50]),.OUT_IBUF(fpgaio_in_int[50]));

	qlIBUF QL_INST_A2F_L_29_3 (.IN_IBUF(fpgaio_in[51]),.OUT_IBUF(fpgaio_in_int[51]));

	qlOBUF QL_INST_F2A_L_30_0 (.IN_OBUF(fpgaio_out_dup_0[52]),.OUT_OBUF(fpgaio_out[52]));

	qlOBUF QL_INST_F2A_L_30_1 (.IN_OBUF(fpgaio_oe_dup_0[52]),.OUT_OBUF(fpgaio_oe[52]));

	qlOBUF QL_INST_F2A_L_30_2 (.IN_OBUF(fpgaio_out_dup_0[53]),.OUT_OBUF(fpgaio_out[53]));

	qlOBUF QL_INST_F2A_L_30_3 (.IN_OBUF(fpgaio_oe_dup_0[53]),.OUT_OBUF(fpgaio_oe[53]));

	qlOBUF QL_INST_F2A_L_30_4 (.IN_OBUF(fpgaio_out_dup_0[54]),.OUT_OBUF(fpgaio_out[54]));

	qlOBUF QL_INST_F2A_L_30_5 (.IN_OBUF(fpgaio_oe_dup_0[54]),.OUT_OBUF(fpgaio_oe[54]));

	qlOBUF QL_INST_F2A_L_30_6 (.IN_OBUF(fpgaio_out_dup_0[55]),.OUT_OBUF(fpgaio_out[55]));

	qlOBUF QL_INST_F2A_L_30_7 (.IN_OBUF(fpgaio_oe_dup_0[55]),.OUT_OBUF(fpgaio_oe[55]));

	qlOBUF QL_INST_F2A_L_30_8 (.IN_OBUF(fpgaio_in_int[13]),.OUT_OBUF(events_o[13]));

	qlIBUF QL_INST_A2F_L_30_0 (.IN_IBUF(fpgaio_in[52]),.OUT_IBUF(fpgaio_in_int[52]));

	qlIBUF QL_INST_A2F_L_30_1 (.IN_IBUF(fpgaio_in[53]),.OUT_IBUF(fpgaio_in_int[53]));

	qlIBUF QL_INST_A2F_L_30_2 (.IN_IBUF(fpgaio_in[54]),.OUT_IBUF(fpgaio_in_int[54]));

	qlIBUF QL_INST_A2F_L_30_3 (.IN_IBUF(fpgaio_in[55]),.OUT_IBUF(fpgaio_in_int[55]));

	qlOBUF QL_INST_F2A_L_31_0 (.IN_OBUF(fpgaio_out_dup_0[56]),.OUT_OBUF(fpgaio_out[56]));

	qlOBUF QL_INST_F2A_L_31_1 (.IN_OBUF(fpgaio_oe_dup_0[56]),.OUT_OBUF(fpgaio_oe[56]));

	qlOBUF QL_INST_F2A_L_31_2 (.IN_OBUF(fpgaio_out_dup_0[57]),.OUT_OBUF(fpgaio_out[57]));

	qlOBUF QL_INST_F2A_L_31_3 (.IN_OBUF(fpgaio_oe_dup_0[57]),.OUT_OBUF(fpgaio_oe[57]));

	qlOBUF QL_INST_F2A_L_31_4 (.IN_OBUF(fpgaio_out_dup_0[58]),.OUT_OBUF(fpgaio_out[58]));

	qlOBUF QL_INST_F2A_L_31_5 (.IN_OBUF(fpgaio_oe_dup_0[58]),.OUT_OBUF(fpgaio_oe[58]));

	qlOBUF QL_INST_F2A_L_31_6 (.IN_OBUF(fpgaio_out_dup_0[59]),.OUT_OBUF(fpgaio_out[59]));

	qlOBUF QL_INST_F2A_L_31_7 (.IN_OBUF(fpgaio_oe_dup_0[59]),.OUT_OBUF(fpgaio_oe[59]));

	qlOBUF QL_INST_F2A_L_31_8 (.IN_OBUF(fpgaio_in_int[14]),.OUT_OBUF(events_o[14]));

	qlIBUF QL_INST_A2F_L_31_0 (.IN_IBUF(fpgaio_in[56]),.OUT_IBUF(fpgaio_in_int[56]));

	qlIBUF QL_INST_A2F_L_31_1 (.IN_IBUF(fpgaio_in[57]),.OUT_IBUF(fpgaio_in_int[57]));

	qlIBUF QL_INST_A2F_L_31_2 (.IN_IBUF(fpgaio_in[58]),.OUT_IBUF(fpgaio_in_int[58]));

	qlIBUF QL_INST_A2F_L_31_3 (.IN_IBUF(fpgaio_in[59]),.OUT_IBUF(fpgaio_in_int[59]));

	qlOBUF QL_INST_F2A_L_32_0 (.IN_OBUF(fpgaio_out_dup_0[60]),.OUT_OBUF(fpgaio_out[60]));

	qlOBUF QL_INST_F2A_L_32_1 (.IN_OBUF(fpgaio_oe_dup_0[60]),.OUT_OBUF(fpgaio_oe[60]));

	qlOBUF QL_INST_F2A_L_32_2 (.IN_OBUF(fpgaio_out_dup_0[61]),.OUT_OBUF(fpgaio_out[61]));

	qlOBUF QL_INST_F2A_L_32_3 (.IN_OBUF(fpgaio_oe_dup_0[61]),.OUT_OBUF(fpgaio_oe[61]));

	qlOBUF QL_INST_F2A_L_32_4 (.IN_OBUF(fpgaio_out_dup_0[62]),.OUT_OBUF(fpgaio_out[62]));

	qlOBUF QL_INST_F2A_L_32_5 (.IN_OBUF(fpgaio_oe_dup_0[62]),.OUT_OBUF(fpgaio_oe[62]));

	qlOBUF QL_INST_F2A_L_32_6 (.IN_OBUF(fpgaio_out_dup_0[63]),.OUT_OBUF(fpgaio_out[63]));

	qlOBUF QL_INST_F2A_L_32_7 (.IN_OBUF(fpgaio_oe_dup_0[63]),.OUT_OBUF(fpgaio_oe[63]));

	qlOBUF QL_INST_F2A_L_32_8 (.IN_OBUF(fpgaio_in_int[15]),.OUT_OBUF(events_o[15]));

	qlIBUF QL_INST_A2F_L_32_0 (.IN_IBUF(fpgaio_in[60]),.OUT_IBUF(fpgaio_in_int[60]));

	qlIBUF QL_INST_A2F_L_32_1 (.IN_IBUF(fpgaio_in[61]),.OUT_IBUF(fpgaio_in_int[61]));

	qlIBUF QL_INST_A2F_L_32_2 (.IN_IBUF(fpgaio_in[62]),.OUT_IBUF(fpgaio_in_int[62]));

	qlIBUF QL_INST_A2F_L_32_3 (.IN_IBUF(fpgaio_in[63]),.OUT_IBUF(fpgaio_in_int[63]));

endmodule

